ELF               �   4 �     4    (        4  4       �   �             �                                     � �          � �      Z  @          �� ��       �           /usr/lib/ld.so.1       �   �           d   �   �   �       >   s                       �   �           �           =                   �   h       �       <       �   �   �           4   �   ^   9          v   �   y   B   u   �                      �   r   �   A   .       +   ]   G       [   �   '       �       �   �   �   H   l   Y   �   �   �   m       C   �       �   -      1   ~   �   x          �   �   k   T   F           w       �   }   W   �           3   X   �   5       O   \   e   �   �   �                   �   _   �   �       R   P      �   i       b   �   o   �   |       �               �                   f                                                                                                                                                                   !               "                                   2                                   *                                           7       8                                   E       L   Q   ;   (       V           ,   S                                          M   g           $               q   J   j       `       n   N       K   6           )   0       c               /              @   z               t       I   �   a   &               {   Z       U   �   p   %   #               �           �       :                  ?   �   D                      �            �                                 �                      8           �           GH      	     GT      
     G`           x`           �           �           ��           ��           �p           �h                                                                                              4�         �        A�   (      ��   �     # �  "     2 �   t     9 h�   �     D FL   x"     I '�   d     [ ��  �     f mp  X     r 4�   "     z 9p   �     � �x        � ��        � �L         � .�   d     � �p          � R@        �    "     � �D  	�     � =�   �     � o�  X     � �  @!     � ��   �     � 4�   l     8�   �     �        - լ   �    C (   d    P A�   ("    Y E�   �"    _ w8      n D�   �    y B8   h"     A�   4"    � �@         � �L         � #@   H    � 1�  �    � .�      � $   �    �     "    � E�  @    � Dd   �"    � *�  �    �        � �|         � F�   �"    � 8$   �    	 >  4     �l  �"     ��  �    . &<   �    ;         A ,�  �    O ��  �    W GH     	  ] �p  �"    b �l  �    h D�   �"    n �   "    s ��         x �      � 6<   �    � ��         � A�   0"    � 'P   d    � D\   "    � ��  �    � c�  0    � @�  4    � �D  	�"    � �  "    � 3�   �    � �x  `"    � ]p         6�   �     ��         \8  �    ! @D   `    4 �d         ; �  @    A #�   D    P D\       Z #�   D    h �  �    o ep       { W`      � :8  H    � 0�   �    � r   X    � ��  �"    � %l   �    � FL   x    � J@       � �X         � �h   X    � B    "    � B         �l  �"     ��   !     �H        tx  X    " H        . B�  �"    5 �l  �    ; B�  �    D ��         I Zh      V ��         ] E�   �    e 4�  �    q �f        x �        � 4�   �    � B8   h    � A�   4    � L@       � ��   �    � �        � G`       � 4(   d    � ��         � Dd   �     ��  �"     (|  T     F�   �     5�   �    ' H  �    , ��       / &�   h    @ ��         E N\  �    P �p  �    W �       ^ D�   �    f 4  x    n N@       { GT     
  � %   d    �     �"    � �x  `    � $�   d    � A�   0    � �  X    � ��         � 7|   �    � �  �"    �     �    � ��   �"   __matherr __sqrt __isnormal __cos _SVID_libm_err _start naf_puiss2 nint i_compl_pdivdoubl naf_iniwin _TBL_cos_hi matherr i_compl_log10 __huge_val _environ _end i_compl_div .stret8 _TBL_log2_lo copysign __expm1 naf_cleannaf _TBL_cos_lo _iob g_NAFVariable i_compl_sub i_compl_log _GLOBAL_OFFSET_TABLE_ cree_list_fenetre_naf i_compl_conj isnormal irint _TBL_ipio2_inf naf_prtabs ilogb isinf atexit exit i_compl_cmplx i_compl_pow i_compl_pow2d i_compl_add log naf_smoy aint i_compl_div2d __copysign malloc rint i_compl_tanh naf_initnaf_notab pow naf_correction i_compl_pmul __log i_compl_div4d __atan2 _init sinh __pow anint fabs .mul __rem_pio2 i_compl_cosh .rem issubnormal i_compl_pmuldoubl signbit __atan naf_four1 naf_mftnaf expm1 sqrt i_compl_exp hypot _TBL_log_hi i_compl_sinh _DYNAMIC naf_inifre naf_cleannaf_notab printf __iob i_compl_module __signbit i_compl_angle __cosh _TBL_log_lo _TBL_atan_hi naf_initnaf i_compl_powreel _TBL_sin_hi atan2 i_compl_mul __nint _TBL_exp2_hi _exit delete_list_fenetre_naf iszero __iszero exp environ errno _TBL_sin_lo __cg89_used scalbn __exp __scalbn free _TBL_atan_lo _write __irint __rem_pio2m _edata _PROCEDURE_LINKAGE_TABLE_ i_compl_cos __ilogb __isinf _TBL_exp2_lo concat_list_fenetre_naf _etext _lib_version i_compl_psub fflush __aint atan i_compl_pdiv __rint i_compl_sin main pi i_compl_muldoubl .div naf_tessol __sinh __fabs __anint __k_sin _TBL_log2_hi _fini i_compl_paddconst sin __hypot i_compl_padd __issubnormal __k_cos fprintf i_compl_tan cosh __sin cos libc.so.1 SISCD_2.3 libc.so.1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �       zt�      �     ��  '     �  k     �x  &     �@  =     �L  >     �X  y     �d  j     �p  *     �|  H     ��  W     ��  �     ��  �     ��  �     ��  Z     ��  �     ��  �    �  ��@��D�, ���@'  ��$���#� �� � � @ ��     �@ ���#T@ JL   � � � � @     @ ��   @ ��   ?��� ch��  	�#�'��  �a��@ �`��@  ����"� �"�  ���h  � ��#  �#   ��cp  ����#� �#�� 
#  ��$`����'  ��$��)  ��%! +  ��%`�-  ��%��/  ��%��1  ��& �� 5  ��&���?�9  ��' �;  �a  ��" �  ��"`��   ��"ਘ   ��#`�  ���p!  � ��$  �$ #  ��cp%  ����$� �$�'  ���p)  � ��%  �% +  ��%`�� /  ��%��1  ��#x3  �`��&@ �&`5  ��&��@ �   �'����������    � l   ;  ��c�  �!��  � ������������V�#�h��h�#�h��h@ 7f     ��#���	X�;�p�����  �!��  � ���\�#�x��x�#�x��x@ 7U     ��c���	B  ������@��p���H����*�  ��`Ğ@�#� �#�!  ��#�  �!��  � ������������R�#�h��h�#�h��h@ 9   #  ��c���	T�;�p�����  �!��  � ���X�#�x��x�#�x��x@ 9   %  ������	\'  ��㘅��@��p���D����- -  ���Į��%��%����� �'��������@���   �      �`��@ �`@ 8   7  ����� ����	��#�h��h�#�h��h� @ �     �� `  ��`�@ ��   � �'��� D   ��h����/`  ������	�� ���"  ���" ���" �" @  V   � ��x����,�)  �� �� �@ �`�"  �`�" �`�" �" @  V   �#�\����.�9  �� �� �  � �#�`�#�d����*�  ��༞��� ������+   ��༞����� ��  �� h� @ �^   ������'�����#  ��`��� ���   �    @ �   �  �    � �����  ?��� c����'�D�'�H�'�L�'�P�'�T��D��H�"  �" ��D��P�# �# �����  ?��� c����'�D��D���� ����D�� ��@ ,�   �    �����  ?��� c����'�D��D���� ����D�� ��@ -�   �    �����  ?��� c����'�D�'�H�����H������D���� �����@�#�`��`�#�`��`��H�� ����D�� ����F�#�d��d�#�d��d���   ����    � @ ��   ?��� c����'�D�'�H��D��H�@ �`�  � ���L�%  �% ��D��H�����������P�%��%������  ?��� c����'�D�'�H��D��H�@ �`�  � ���T�&  �& ��D��H�����������X�&��&������  ?��� c����'�D�'�H�����H� � ��D�`�`���\��H�@ �`��D�� �����@�����#�`��`�#�`��`��D������H�  � ���H��H�`�`��D�� ����	J��F�#�d��d�#�d��d��I   ����    � @ ��   ?��� c����'�D�'�H��D�� ���?����H�`�`��D�������P��H�� ��������T������D�%  �% ��D�`�`��H�� �����\��H���������	^��Z��D�& �& �����  ?��� c����'�D�'�H�'�L��L�@ �`��D��H���D�?����L������D��H���H�?������    � @ �J   ?��� c����'�D�'�H��D��H�  � �� �����L�&� �&���D��H�  � �`�`���P�'`�'`�����  ?��� c����'�D�'�H��D��H�� ���@ �`�����"@ �"`��D��H�  � ���������"��"������  ?��� c����'�D�����D���� ���� ��#�`��`�#�`��`��D�� �����   ����    � @ ��   ?��� c����'�D�'�H��H�@ �`�?��#  ��c���聨
�      	�    �    %   �����'����H� � �'���'��-  ���������
�      	�    �    /   ��� �'������������      �    � 1   ��H�`�`��H�� ����	��?�����������P7  ��㨩��N��H� � ���T�?����D�@ �`�����	Z��D� � ��\��𽧉��?����D�`�`������D��D�� ���������	���D�"��"�� /   ��H� � ��H�@ �`��	��?����������	R  ��㨭�P��H�  � ��	V�?����D�`�`������\��D�� �����Z�����	��?����D�� �������	F��D� � �����𕢉���D�%`�%`��D����%� �%������  ?��� c����'�D�'�H�'�L�'�P�'�T�'�X��L��P5  ��������      	�    �    �� :�� ;�� ��� 0�� 1��T��X7  ��㰁�
�      	�    �    �� 8�� 9�� ��� 4�� 5����      �    �     ��L��P��T��X������ 6�� 7�� >�� ?���^9  ��#���B��T��X��	F�� (�� )��D��H���^�����?����D��H�� ���	��?���    ��T��X��L��P���н� .�� /�� >�� ?���^;  ��c���R��L��P��	V��  �� !��D��H�����?����D��H�� ���	^��	��?������    � @ ��   ?��� c����'�D�'�H�'�L�'�P�'�T�'�X��T��X  ��#�����      	�    �    �� :�� ;�� ��� (�� )��\��`  ��c���
�      	�    �    �� 8�� 9�� ��� ,�� -����      �    � &   ��T��X��\��`���н� .�� /�� >�� ?���^  ���ȭ�R��\��`��	V��  �� !��D��H���^��L��P���D�����?����L��P��	^��D��H��ʙ�	��?��� $   ��\��`��T��X���н� .�� /�� >�� ?���^  ���ȭ�R��T��X��	V��  �� !��L��P���^��D��H��B�����?����D��H��	^��L��P���ș�	��?������    � @ �~   ?��� cp���'�D�'�H�����D�@ �`�#  �`�# �`�# �# �����H��n   ����    � @ �e   ?��� cX���'�D�'�H�'�L�'�P�'�T)  ��#й� .�� /+  ��cص� 0�� 1��T�� �    �    � d   ��T�� �    � '   ��T�  �'�T  ��#���D��H��L��P����#�@�;�`�;�h�;�p�;�x�;�����      ��`��h��p��x�������  � �&� � �&�� �&��&��������    ��D��H��L��P��T��`�    �    �� :�� ;���V�� <�� =��	X��ҽ�  �� !�� :�� ;���X�� <�� =��	V��B�� &�� '�� >�� ?�7`�� �    �    �� 6�� 7��	V�� 8�� 9���X���Ƚ� ,�� -��X���N�� >�� ?�    �    ���   �?���?������    � @ ��   ?��� cX���'�D�'�H�'�L��`��D�� ���"  ���" ���" �" ���   �;�p��p��t��H@ ,
   �?����`��D�  � �"  � �" � �" �" ���   ��H��	@�?�����@ 3   ������@�?�����@ 4�   �����	@�?�����    � @ ��   ?��� cp���'�D�'�H���7  ������ ���&� ���&����&��&���H�� 
�    �    � W   ��H�� �    �    ��H�  �'�H  �����?��!  ��#��?�ؐ����D���   � 
   ��D�@ �`�?����D�����?����H�'���������    �    �����ص��\�����н��@�����?�������Љ�	F�����ؑ�	J��D�?������?������6��'������� �    �    �����؝��P�����Х��T�����?����е�X��ع�	Z�?������?���    �    ���   ����    � @ �6   ?��� c����'�D��D�� ��@ 2�   �?����D���� ��@ 2v   ��轧�@�?����D���� ��@ 4I   ��腠�@�?������    � @ �   ?��� c����'�D�'�H��D��H�@ �`�  � �����"  �" ��D��H�������������"��"������  ?��� c����'�D�'�H��H�  � ��D�@ �`�����?����H������D� � ����?������    � @ ��   ?��� c����'�D��D���� ��@ -�   �;�`��D�� ��@ 2    ��`��	X�?����D���� ��@ .G   �;�`��D�� ��@ 3�   �� ���`��	Z�?������    � @ ��   ?��� c����'�D��D���� ��@ -�   �;�`��D�� ��@ 3�   ��`��	\�?����D���� ��@ .   �;�`��D�� ��@ 1�   ��`��	^�?������    � @ ��   ?��� c����'�D��D���� ��@ 1�   �;�`��D�� ��@ -�   ��`��	B�?����D���� ��@ 3�   �;�`��D�� ��@ -�   ��`��	D�?������    � @ �g   ?��� c����'�D��D���� ��@ 1�   �;�`��D�� ��@ -�   ��`��	F�?����D���� ��@ 3z   �;�`��D�� ��@ -N   ��`��	H�?������    � @ �?   ?��� cp���'�D��D�@ �`���J�?����D�������N�?�����@ -4   �;�`���@ 1z   ��`��R�?�����@ 3P   ��؁�	��?�����@ -�   ��؁�	��?������    � @ �   ?��� cp���'�D��D�� �����Z�?����D� � ���^�?�����@ -
   �;�`���@ 1P   ��`��B�?�����@ -z   ��؁�	��?�����@ 3    ��؁�	��?������    � @ ��   ?��� cx���'�D��`��D�@ �`�"  �`�" �`�" �" ���   �;�p��p��t@ 2B   �?���`��D�� ���"  ���" ���" �" ���   �?������    � @ ��   ?��� cp���'�D  ��  @ 2&   �?���`��D�  � �"  � �" � �" �" ��s   �;�p��p��t@ 2   ��聠	��?���`��D�  � �"  � �" � �" �" ��p   ��聠	��?������    � @ ��   ?��� c���5  ���7  ����&� �&�9  �!��  � ��P  � ��  � ��	�  �`��"@ �"`  ������  ����� ����	Z  � ��  � ��	�  �`��#@ �#`  �� �� �* @ �e   �'�����!  ��$ ������ �    � 	     �� �@ �Q   � @ �H     �� �� �* @ �N   �'�����'  ��$������ �    � 	     �� �@ �:   � @ �1     �� ��   ��`��`@ �8   �* @ �2   � �� �    � 	     �� �@ �"   � @ �     �� �� �* @ �   �'�����-  ��%������� �    � 	     �� �@ �   � @ �   �'���    ����. 5  �����&�7  �������/ �@����`�'��  ��������� ���   �      �� �� �* @ ��   �'�����  ��#����� �    � 	     ��!@ ��   � @ ��     �� �� �* @ ��   �'�����%  ��$������� �    � 	     ��! @ ��   � @ ��     ��!�@    �����  ?��� c���  �� �@ ��     �� �@ ��   )  �� ��  @ ��     �� �@ ��     �� �@ ��     ��!�@ ��     ��! @ &   +  ��%a �����  ?��� c���-  ���/  ����%� �%�1  �!��  � ��@3  �`��@ �`��	�5  ����&� �&�7  ������9  � ��  � ��	J  � ��  � ��	�  �`��"@ �"`  �� ��   ��`��`@ �p   �* @ �j   � �� �    � 	     ��!8@ �Z   � @ �Q     �� �� �* @ �W   �'�����  ��"������� �    � 	     ��!P@ �C   � @ �:   �'���    ����+`!  �� ��$ #  ��`��`�,��@���� �'��+  ��`��`���������   �      �� �� �* @ �'   �'�����3  ��&a������ �    � 	     ��!h@ �   � @ �
     ��!�@ c   �����  ?��� c���7  ������ @ �     �� �@ �
     ��!�@ �     ��! @ %w   9  ��'! �����  ?��� c8���'�D�'�H�'�L��D  �� ���@�    � 	     ��!�@ ��   �  � �     ��`�?��  �`��@ �`@ 07     ��� ��	��?��@ �     �� �� ���@ 	�     ������  � ��  � ���T����������?��  ��a �� �    �    ����'������'��� W   ����4`���<`�$`�'��)  ��! � �'�D-  ��� �� �������	ށ�\�'��/  ��� ����������č�B�'���������� �    � 
   ������?������'�������J�'������  �����@�    �    ����  �'���    ����������    �    ����'������  ����� �    �    ����  �'���    ����������    �    ����'��� �'�������D����    � P   ������������@ �   �?����H�#�\�#�`��ؒ�Д�Ȗ�����@ �   ������������ � @  �   ����� �    �    � /   �����`�    �    ���������@ K   �� �    �    �  � 7     ������  ��"������?��    �    ��Д�����@ 	�   ����`�'�������D������   �    #  ��a �� �    �    %  ��� �'�������+  ��%a ���@ ��   -  ��� �� ��3   �    � �    � �����  ?��� c����'�D�'�H�'�L/  ��ഀ���    � *   �'�������D�� �    � "   ����.���H� �`�`�;�X����*`��H��
�� ��  ��a����  �� ���X@ ��   ��L���� �'�������D��@���   �    �����  ?��� c����'�D!  �� �� �#�`��`���?��%  ���(� � )  �� (� � ��D��O   �'��-  �����'���    ��D������   ������'������'������`�'�����7  ����������   �    �����D��N   �'��9  �� ��'���    �����D��a   ����`�'������'������`�'�����  ����������   �    �����  ?��� c����'�D�'�H�'�L�'�P�'�T�'�X��L� �#    �`��@ �`@ .�   �?�� �'��� f   ����,   ��พ��� ����D��H����#�`��`�#�`��`@ .�   �?������������      	�    � I   �����𵦉���P����      	�    �    ��L�?��$� ��X����%  -  ��������    �      �� �  ��a���������	��#�`��`�#�`��`@ �   � -   ��L�%� 1  �� ��� �    �      �� �  ��a�������@ �   ����.`  ��พ��� ��  ��a���D��H  �� �@ ��   ������'�����;  ��`��� ���   �    �����  ?��� c0���'�D�'�H�'�L�'�P�'�T��H�" ��D���	�    � 	     ��"$��D@ ��   �>   ��`��T�� ���"  ���" ���" �" ��p��P�� ���"` ���"`���"`�"`����#�@���      ��L�  � �&` � �&`� �&`�&`� �'����L�`�'�������H����    � 4   ��`��Ğ#`�� ���"  ���" ���" �" ��p��P�  � �"` � �"`� �"`�"`����#�@���      ����  � �&� � �&�� �&��&����� �'������'����Ğ��'�������H�� ���   �    ��`��H�,���L� �%`�� ���"  ���" ���" �" ��p��T�  � �"` � �"`� �"`�"`����#�@���      ����  � �$  � �$ � �$ �$ ���-  ���0� � 1  �� 8� � ���   �'����D� ��H@ �=   �'�� �'�������쀦��    � P   ��Ȓ�����   ��H���� �'���'�������H��@
�    � 6   ��`����*���L�@�� ���"  ���" ���" �" ��p����  � �"` � �"`� �"`�"`����#�@��8      ���������/`��L��	�  � �"� � �"�� �"��"�������'�������H������   �    ���`�'�������쀥����   �    ��Ȓ����E   ��H����@�'�������H@ ��   �  ��D��� �'���'�������� 	�    � 6   ��`����*���L� �@ �`�"  �`�" �`�" �" ��p����  � �"` � �"`� �"`�"`����#�@���      ���������/`��L��	�  � �"� � �"�� �"��"�������'������������   �    �����  ?��� b����'�D�'�H�'�L�'�P�'���'���'���'��  �� �� �* @ �y   �'������� �    � 	     ��"8@ �h   � @ �_     �� ��   ��`��`@ �f   �* @ �`   � �� �    � 	     ��"P@ �P   � @ �G     �� �� �* @ �M   �'������� �    � 	     ��"h@ �<   � @ �3   �'�|�    ��|�-�����&@5  �������.��@��|� �'�|  ��`��`��|���
���   �      �� �� �* @ �!   �'������� �    � 	     ��"�@ �   � @ �     �� �� �* @ �   �'������� �    � 	     ��"�@ ��   � @ ��     ������!  � ��  � ���H�?���'��#  ��`��'���    %  ���@� � )  �� @� � ������   ������'������'�|���� �'�����5  ������@���   �    ���  ���@� 
�   �� H� � ��{   � �'����   ��`����  � �"� � �"�� �"��"�����-�  ��พ��� ��1  � ��  � �����#�p��p�#�p��p��x�#�@��C      ����  � �&� � �&�� �&��&��������, %  �������� ���#� ���#����#��#�1  �� ��� �    � �   �������@ �`�"� �`�"��`�"��"�  � ��  � ��襣�P  ����� �������#������#���������#�@��      ����  � �#` � �#`� �#`�#`� ����#�@��&      ��p�  � �"` � �"`� �"`�"`��`����� ���"  ���" ���" �" ����#�@��      ����  � �$  � �$ � �$ �$ ��p����� ���"� ���"����"��"�  �`��@ �`����#�@���      ��`�  � �"` � �"`� �"`�"`� 	����#�@���      ����  � �$  � �$ � �$ �$ ��`����� ���"� ���"����"��"���p����  � �#  � �# � �# �# � @���  �� ���   �'��%  �����'���    ����,�����@������   ����`�'������'�x������'�����3  ��`��� ���   �    � �   �������� ���"� ���"����"��"�  � ��  � ��蹦Z  ����� ������#������#���������#�@��U      ����  � �$` � �$`� �$`�$`� ����#�@��t      ��p�  � �"` � �"`� �"`�"`��`����  � �"  � �" � �" �" ����#�@���      ����  � �$  � �$ � �$ �$ ��p����� ���"� ���"����"��"�  �`��@ �`����#�@��      ��`�  � �"` � �"`� �"`�"`� 	����#�@��1      ����  � �$  � �$ � �$ �$ ��`����� ���"� ���"����"��"���p����  � �#  � �# � �# �# � @���  �� ���g   �'���    ����,�)  �� Ī �'�x����-����� �@ �`��x�� ����B�&� �&�������'�����  �� ��� ���   �    ����`�'�����  ��ࠀ����W   �    ���@ �   � �'��� I   ����+`���� ����,�)  �� �� �@ �`�$@ �$`����-�����@����.�  �� �� �@ �`�&� �`�&��`�&��&�� �'���    ����, ���������- ������-�3  ��`��@����.����  � �%� � �%�� �%��%�������'�����#  ��`��� ���   �    ������'�����)  �� �������   �    +  ��`��'�������D��H���   �� �    �    ����� @ ��   ���@ ��   ���@ ��   ���@ ��   �  � �   � �'��� #   ����. ��L������/   ��`��@�� ���&� �&�����+ ��P������,`'  ��༨��  � �$  � �$ � �$ �$ ������'�����9  �� �������   �    � �'��� I   ����*`  ��ธ�
����+`���� �@ �`�#  �# ����,�+  ��`��@����-�����@�� ���%� ���%����%��%�� �'���    ����+`!  �� �� ����,��@����-`���������.`� �� ���%  ���% ���% �% ���� �'�����  ��ࠀ�@���   �    ���� �'�����%  ������@���   �    ����� @ �(   ���@ �%   ���@ �"   ���@ �   � �    � �����  ?��� c���)  �� ��'��+  ��`P�?��-  �������'��1  �� �� �'�� �'����������    � H   ����/`  ��`��@�'���������"� �"������'���������$  �$ ��� �'���������%@ �%`��� �'�� �'�������􀦀�    �    �������'  �' ��ܔ��'���������"� �"���ܞ��'������ �'��������@���   �    ������'�������� ���   �    -  ��%�������  ?��� c@���'�D�'�H�'�L�'�P�'�T�'���'����T�'����Բ& �'����Ԑ �* @ ��   �'������� �    � 	     ��"�@ ��   � @ ��   ��ԑ* @ ��   �'����܀� �    � 	     ��"�@ �x   � @ �o   9  �� ��� �    �      �� �  ��b������L��P@ �t   �?��'����ԕ��?�Ȑ �'���'������'��  �����'�������؀���    � 4   ���+`!  ��!�� �@ �`����� �����L����$� �$����� �'����Ī`�'�����-�1  ��!�� �@ �`����� �����P����&� �&����� �'����ĺ`�'����� �'�������؀�@
���   �    ����" ������@  �   �'������'����Ě �'�������؀���    � /   ����@ �`����� �����T����� ������� �����X���V�#�p��p�#�p��p@ *	   ��ȁ�	����- ��ܮ��%� �%���� �'����Ĳ`�'��������'�������؀�����   �    ���@ ��   ��D��Ԁ�@�    �    ������@    �'����ԕ2`��	�:`������ 	�    �    ����'���    �����Ԣ#��'������'��� `   ��D�� �    �    ��H��D�" ��D�-`��ܒ@@ �   ��D���'������'��� J   ��H�� �    �    ��H��D�" ��Ի/ ��ܒ@��D�*��@@ �   �'�������D� �'��� 1   ��D�  �" ��ԣ, ��ܒ@��D�,��@@ �   ��D� �'����H���@ �   �'�������԰��. ��ܶ��� �����/ ��ܒ �@ �`����      	�    �    ����'���    ����'����䍠��L��P���H���
���L�?��  �� ��� �    �    ���+`��ܢ �@ �`�;�`����;�X����#�h����#�l  �� �  ��b���D��H�����X@ �C   ���@ �=   ����    �����  ?��� c@���'�D�'�H�'�L��H� �'��� �'��� �'���������� �    � g   �������� 	�    � 7   ����*���D� �@ �`�?������,`��D��� � �'���'������-���D� ����.���D� �@ �`�&@ �&`����*`��D��
����+`��D� �`�`�# �# ����,���D�@����%� �%�����.���D� ����'`�'`����2���
�:��'��� 	   �������#@�'�����;��'������� �    � 	   ��������@���   �    ������� �'������`�'��������������   �    � �'�������쀦@�    � �   �����'����L���@ ��   �#�`��`��;  ��`X�����?��  �� `��୥�T�#�`��`�#�`��`@ '�   �?��  ��`h������X������\�?�����@ '�   �?��  ���p�?��  ���x�?��� �'�������쀣@�    � �   ����'����������@�    � e   ��������'������-���D� �`�`�����	B����.���D� �@ �`��ȑ�	F����?������* ��D��	�� ��������L����+ ��D��� � ��ȥ��P���N�?������,`��D���  � �����������-`��D���&  �& ����.`��D��� � ����������/`��D�@�"��"�����*���D�@����� ����B�#� �#�����, ��D�����������F�$��$��������@�'��������������   �    ����?�������Е��L�����؝��P������ȩ�R�?�������Э��X�����ص��\���V�����^�?�������'�������쀦���x   �    ����'�������쀢 	��<   �    �����  ?��� c����'�D�'�H��D�'������� �    �    ��H�#  �    ��H� �#@ ����� �    �    ��H��H�� ���$@ ����=`�'�����������   �    �����  ?��� c����'�D�'�H�'����H�� ���?�� �'�������D����    � #   ����/ ��H� �@ �`�������      �    �    ����*���H� �@ �`�?������'��������'�������D������   �    ����    � �����  ?��� c����'�D�'�H� (�'���'������������    �    1  �� �����.`��H���'  �' ;  ��`���D����" 	�*���H� �#@ �#`������'���������� ���   �    �����  ?��� b����'�D�'�H�'�L�'��%  �����'��  �� �� �* @ �E   �'������� �    � 	     ��#4@ �4   � @ �+   ���)  �� �� � -  ����� � ���   ��x����  � �"� � �"�� �"��"���D�*   ��พ�	�� ��  ����� �������#������#���������#�@��      ����  � �#` � �#`� �#`�#`�����H�� ����L�� ����   ��x����  � �"  � �" � �" �" ��   �;��������  �� �  ��cL��D@ ��   ��D�.�  �� �� ������   9  �� ��� �    � F   ��x��D�/`  ������	�� ���"  ���" ���" �" ��   �;����D�,�  ��༞����� ����D�-   ��༞��� ��@ �   �#�l�#�p��D�-�1  �� �� �@ �`�#�\�#�`��D�.�;  ��`��@� � �#�d�#�h��D�*�  ��พ��� ��  ��ct  �� ����@ ��     �� ��� �    � �   �������@ �`�"� �`�"��`�"��"�  � ��  � )  � ��  � �����#������#���������#�@��      ����  � �%� � �%�� �%��%�� ����#�@��*      ����  � �"` � �"`� �"`�"`��x����� ���"  ���" ���" �" ����#�@��      ����  � �%` � �%`� �%`�%`�������� ���"� ���"����"��"�  �`��@ �`����#�@���      ��x�  � �#  � �# � �# �# � ����#�@���      ����  � �%` � �%`� �%`�%`��x����� ���"� ���"����"��"��������� ���#  ���# ���# �# � @���  �� ���   �'��)  �� ��'������'������������    �    ���������   ���� �'������'��������'������'������ �'����������@���   �    � �   �������@ �`�"� �`�"��`�"��"�  � ��  � %  ����� ������#������#���������#�@��S      ����  � �%  � �% � �% �% � ����#�@��r      ����  � �"` � �"`� �"`�"`��x����  � �"  � �" � �" �" ����#�@���      ����  � �%` � �%`� �%`�%`�������� ���"� ���"����"��"�  �`��@ �`����#�@��      ��x�  � �#  � �# � �# �# � ����#�@��/      ����  � �%` � �%`� �%`�%`��x����� ���"� ���"����"��"��������� ���#  ���# ���# �# � @���  �� ���e   )  �� ���D�-`/  ��ะ��  � ��
Z      �    � (   �'����������@�    �    ����.�;  ��`Đ@�'������*`�����
�  � ����@ �`����#@ �#`������'���������� ���   �    � '   �'������������    �    ����- -  ���Į��'������. ������� �����B����  � �����'  �' ����`�'���������� 	���   �    ���@ ��   �����  ?��� bX���'�D�'�H�'�L�'�P�'�T�'�X�'���'�d  �����'�X  �� �� �* @ ��   �'�d��d�� �    � 	     ��#�@ ��   � @ ��     �� �� �* @ ��   �'����܀� �    � 	     ��#�@ ��   � @ ��   � �'��� "   ����+�  ��พ��� ������,`��ܘ ��D��H@ �   �� �    �    ��d@ ��   ���@ ��   �  ��   ������'�����+  ��`��� ���   �    -  �������'�����. ��ܐ 5  ����� � 9  �� �� � ��   ���*   ������	��D��H�"� �"�� �'��� �   ����'��� u   � �'����������@�    � i   ����,�+  ��`��@����-�� ����#�@��/      ����  � �&` � �&`� �&`�&`� �������*�  �� �� ����+��@�@ �`�"` �`�"`�`�"`�"`����#�@��d      ��x�  � �%� � �%�� �%��%�� �������/ ��ܖ��� ���"` ���"`���"`�"`����#�@��H      ��H�  � �$� � �$�� �$��$����. 5  ����������.�� ��H���   ����`�'���������� 	���   �    ������'�����  �� �������   �    ����`�'�����!  �� ������z   �    ���,`'  ���������- � -  ����� � 1  �� �� � ��v   5  �����?�����9  �� �� �   �� �� � ��h   � �'���������� �    � B   ���,�)  �� �� ����-`� ����#�@��      ��x�  � �&  � �& � �& �& � �������*���ܚ �@ �`�"` �`�"`�`�"`�"`����#�@���      ��H�  � �%` � �%`� �%`�%`��Ȓ�H��   ������'��������������   �    ��x����@ �`�"  �`�" �`�" �" ��%   �;��������@ #i   �?��  ��ഀ���    �    ����#�\�#�`  �� �  ��c�������@ �S   � �'������������    �    ���-`/  ����������. � �����   ������'��������������   �    �����L��P��������#�x��x�#�x��x��T��X��������#�|��|�#�|��|���   ���  ����� 
�   �� �� � ��   � �'���������� �    �V   ��x����� ���"� ���"����"��"�����.   ��พ��� ��5  ����� �������#������#���������#�@��      ��h�  � �'  � �' � �' �' ��x���+�#  ��`��@����,����@ �`�"  �`�" �`�" �" �������� ���"` ���"`���"`�"`����#�@���      ��x�  � �#` � �#`� �#`�#`����-   �� �� ��x��   -  ��������    � F   ��x����-�3  ��`��@�� ���"  ���" ���" �" ��X   �;������+   ��༞����� ������+�  ��༞��� ��@ Z   �#�l�#�p����,`'  ��༨��  � �#�\�#�`����-�1  �� �� �`�`�#�d�#�h����.�  ��พ��� ��  ��c�  �� ����@ �j   ;  ��`���`�    � �   �����h�  � �"� � �"�� �"��"�  � ��  � %  ����� �������#������#���������#�@���      ����  � �%  � �% � �% �% � ����#�@���      ����  � �"` � �"`� �"`�"`��x��x�  � �"  � �" � �" �" ����#�@��T      ����  � �%` � �%`� �%`�%`�����h�� ���"� ���"����"��"�  �`��@ �`����#�@��      ��x�  � �#  � �# � �# �# � ����#�@��      ����  � �%` � �%`� �%`�%`��x����� ���"� ���"����"��"��������� ���#  ���# ���# �# � @��d  �� ����   �'��)  �� ��'�`��d�'�\�����X����    �    ��`��\��   ��� �'����`�'�P��`���'�`��\�'�T��\� �'�\�����X��@���   �    � �   �����h�@ �`�"� �`�"��`�"��"�  � ��  � %  ����� ������#������#���������#�@��"      ����  � �%  � �% � �% �% � ����#�@��A      ����  � �"` � �"`� �"`�"`��x��x�  � �"  � �" � �" �" ����#�@��      ����  � �%` � �%`� �%`�%`�����h�� ���"� ���"����"��"�  �`��@ �`����#�@���      ��x�  � �#  � �# � �# �# � ����#�@���      ����  � �%` � �%`� �%`�%`��x����� ���"� ���"����"��"��������� ���#  ���# ���# �# � @��d  �� ���4   )  �� ���D��H��
B      �    � (   �'�������X��@�    �    ���-�3  ��`Ĵ@�'�T���.���d�@�  � ��T�@ �`����"@ �"`�����'�������X������   �    � '   �'�������X��@�    �    ���, %  ���Ħ��'�T���- ��d���� �����J��T�  � �����&  �& ���`�'�������X������   �    ���� �'����������@���   �    ��d@ �   ���@ �   � �    � �����  ?��� bp���'�D�'�H�'�L�'�P�'�T���  ����� 
�   �� �� � ��C   ��D��H  ����� ����	��?����L��P!  � ��  � ��	��?�x%  ����� ���'���'��%  ������'  ����� �����\)  � ��  � ���Z�?����h����@ �`�"� �`�"��`�"��"����������������x��ʙ�	F�#�x��x�#�x��x����#�@���      ����  � �&� � �&�� �&��&���h����  � �"� � �"�� �"��"������x����������T�#�x��x�#�x��x����#�@���      ����  � �%` � �%`� �%`�%`��h����� ���"� ���"����"��"������x����������\�#�x��x�#�x��x����#�@��      ����  � �#  � �# � �# �# �������  � �"  � �" � �" �" ����#�@���      ����  � �'` � �'`� �'`�'`��Ȟ���� ���"  ���" ���" �" ����#�@��      ����  � �"` � �"`� �"`�"`� ����#�@���      ��h�  � �&� � �&�� �&��&�� ��x����  � �"` � �"`� �"`�"`����#�@��<      ��T�  � �%` � �%`� �%`�%`5  ����� ��7  ���� �����@�?������������9  �� ����H�?�������x����������P�?�����������T��������?�����@ �   ;  ��`���
�      	�    � <     �� ��#�\  �!  ��`  ����� ��  �`��@ �`@ ~�     �!  ��`H��D��H��L��P@ ~v   ����#�\�#�`  �!  ��`X������@ ~k   ����#�\�#�`  �!  ��`p�����x@ ~`     �!  ��`����@ ~Y   �    ����� ������	��?�������T���   �����  ?��� c����'�D�'�H���  ��p  ��h��D��H@ L   ����    �����  ?��� c����'�D�'�H��������D��H  ��p  � h@     ����    �����  ?��� b����'�D�'�H�'�L�'�P�'�T�'�X�'�x  �� �� �* @ ~   �'�x��x�� �    � 	     �� �@ }�   � @ }�   ��D��H!  � ��  � ��	��?�����%  ���Ȓ � )  �� Ж � ��   -  �����'�|���/  ����� ����	F�?�����1  � ��  � ��	J�?��������@ �`�"� �`�"��`�"��"���� ��#������#���������#�@��a      ��p�  � �#  � �# � �# �# � ����#�@��      ����  � �%` � �%`� �%`�%`�������� ���"� ���"����"��"���蝠 ��#������#���������#�@��4      ��p�  � �#  � �# � �# �# � ����#�@��S      ����  � �%` � �%`� �%`�%`��p����� ���"  ���" ���" �" �������  � �"` � �"`� �"`�"`����#�@���      ����  � �%` � �%`� �%`�%`�������� ���&� ���&����&��&��#�\��p����� ���#` ���#`���#`�#`� @��x  ����  ��!�  �� �@ i   )  �� ���|����	��?�������|�����x@ �   ��P����%@ �%`��T����&  �& ��p����  � �"  � �" � �" �" ���   ��X�#� �#��������@ �`�$  �`�$ �`�$ �$ �#�\/  ����� ���;�`3  �`��@ �`�;�h��p����@ �`�#` �`�#`�`�#`�#`� @��x  ����  ��!�  �� �@  2   �����|�����x@ t   �������#�@���      ��p�  � �"� � �"�� �"��"�� 
�������� ���"` ���"`���"`�"`����#�@��      � � ���V��L�&@ �&`��x@ |�   �����  ?��� b؝��'�D�'�H�'�L�'�P�'�T�'�X�'����H�* @ |�   �'����Ā� �    � 	     �� �@ |�   � @ |�   ��H�&���D��@�    �      �!  ��`���D@ |�   �   ��`��\�@ �`�"  �`�" �`�" �" ��p��X�� ���"` ���"`���"`�"`����#�@��      ����  � �%` � �%`� �%`�%`� �'�������H����    � 5   ��`����/`��Ė�	�"��  � �"  � �" � �" �" ��p��X�  � �"` � �"`� �"`�"`����#�@��      ����.���Ē@�  � �"` � �"`� �"`�"`������'�������H�� ���   �    �'�������H����    � V   ��p����- ��P���� ���"  ���" ���" �" �������/ ��Ė��� ���"` ���"`���"`�"`����#�@��N      ��`�  � �"� � �"�� �"��"��������h��	^��`��\����. ��T���� �����D�#������#���������#�@��      ����/`��L��	�  � �"� � �"�� �"��"�������'�������H������   �    ��`��H�-`��İ��& �@ �`�"  �`�" �`�" �" ��p��\�� ���"` ���"`���"`�"`����#�@��A      ����  � �$� � �$�� �$��$����1  �� ؒ � 5  ����� � ��\   �'����D� ��H@ {�   �'��� �'��������@�    � �   ��Ȓ����   ��H�����	�'���'�������H����    � x   �������+`��Ģ �@ �`�"  �`�" �`�" �" �������� ���"` ���"`���"`�"`����#�@��      ����  � �"` � �"`� �"`�"`��p���������,`��P���  � �"  � �" � �" �" ����#�@��      ��`�  � �"� � �"�� �"��"����������#����Б���h��	J��`��H���������- ��T���� �����P�#������#����԰���#�@���      �������@�.���L�@�  � �"` � �"`� �"`�"`������'�������H�� ���   �    �����'�����������t   �    ��Ȓ����w   ��H������'�������H@ {   �  ��D� �`�'���'�������쀦��    � x   �������/`��Ė�	�� ���"  ���" ���" �" �������� ���"` ���"`���"`�"`����#�@��      ����  � �"` � �"`� �"`�"`��p���������+ ��P���  � �"  � �" � �" �" ����#�@���      ��`�  � �"� � �"�� �"��"�������� �#����Щ���h��	V��`��T�������@�+ ��T���� ����	Z�#������#����Ԟ���#�@��0      ������� �,���L� �  � �%` � �%`� �%`�%`������'�������쀦����   �    ���@ z   �����  ?��� c8���'�D�'�H�'�L�'�P�'�T�'�X;  ��'`�  � ��  � ��T��X����      	�    �    ��T��X�'���'���      ����� ���?������?����L��P@ �   �����
�      �    �    ��`����    �    ��d  ��`�@ zD   �'����D��H��L��P����?����D��H�?�������    �?�������蝢���#�h��h�#�h��h@ �   �����
�      �    � �   ����?��������   �?�������ح����?����`�� �    �    �����蹦��#�h��h�#�h��h@ `   �#�\�#�`��d  ��`�������@ z   ��d  ��a������@ y�   ���@ M   +  �`��@ �`��
�      �    �     � /  ��%���`�� �    �    ��d  ��a4@ y�   ��d  ��aX@ y�   ��d  ��at@ y�   ��\����&@ �&`� �   �����������Ѝ��D��ȍ����?������?����������J�?������ �'�������`�    � !   �   ��"���`�� �    �    ��d  ��a�@ y�   ��d  ��a�@ y�   ��d  ��a�@ y�   ��\��D��H�#@ �#`� Z   ��d   ��\����$@ �$`�����𥣈P�#�h��h�#�h��h��T   �;�p��������#�x��x�#�x��x��J   ��p��	Z)  �� 聨
�      �    �    � -  ��%����`����    � -   ��\�� ��  ��b��d���@ yd   1  �� ��� �    �    ��d  ��b,@ yX   3  ��`��� �    �    ��d  ��b<@ yL   ��\�� ��  ��bL��L��P��d@ yB   �����  ?��� b����'�D�'�H�'�L�'�P�'�T�'�X5  �����?��7  �����?��  �`��@ �`@ .   ��T��X����      	�    �      �`��@ �`@    �?���    ��T��X�?������?����d����    �    ��h  ��b`@ y	   ��L��P�'���'���'���'��  ��# ���D��H�?��������   �?����������?�������𝢈L�?��������   �?��������   �?�������`�� 
   �    ������d�    � D   ������d�    �    � +  ��%`���d�� �    �    ��h  ��b�@ x�   � *   �����L��P��
�      �    �    � 1  ��& ���d�� �    �    ��h  ��b�@ x�   �    � 7  ��&���d�� �    �    ��h  ��b�@ x�   ����?����   ��������
�      �    �    ��������
�      �    � *   ������'����������
�      �    �    ����?������?���    ����?������?������������?�������𕡈H�?�������   �?�������   �?����z   �����ȡ���?�������������?�����������-  ������	^��������	B��	��#������#�����@ �   �?����d����    � 7   ���@ C   1  �� ���
D      �    �    ���@ 7   ��荡���#�t�#�x����#�\�#�`����#�d�#�h����#�l�#�p��h  ��b�������@ x    �    ����#�\�#�`����#�d�#�h����#�l�#�p��h  ��c������@ x   ���@ _   %  ��� ��
�      	�    �    ���@ S   �?�x�    '  ��� �?�x����������#������#�����@ D   )  � ��  � ���R��x��	V��
�      	�    �    � -  ��%����d����    �    ��h  ��c4@ w�   ����?���   ���@ !   5  ��� ��
�      	�    �    ���@    �?�p�    7  ��� �?�p9  � ��  � ��p��	^�����
�      	�    �    �   ��" ���d��`�    �    ��h  ��cP@ w�   ����?��� �   ���@ �     ��! ����      	�    �    ���@ �   �?�h�      ��a �?�h��h��������#������#�����@ �   ��蕢�@�����
�      �    � ,   ��d����    �    ��h  ��cd@ wh   !  ��! �������      	�    �    ����?�`�    )  ��! �?�`��`�����	��#������#�����@ Q   ��豦	@�?��� �   +  ��`����	Z������������	B��������ƹ�	��?�����@ �   -  ��� ����      	�    �    ���@ �   �?�`�    /  ��� �?�`���@ x   1  � ��  � ��`���P��
�      	�    �    ��d��`�    �    ��h  ��c�@ w   ����?��� ?   ���@ Y   �?��9  �� ������
�      �    �    ����?������?�������ر�V�?��������   �?�������𽦈\�?��������   �?���    ����?������?�������؅����?��������   �?����������?��������   �?��������'�����   ��\����$� �$���`����%� �%���d����    � U   ��`�� ���#�\�#�`��\�� ��  ��c������h@ v�   ��h  ��c����@ v�   �����ȝ����#������#�����@ �   �;������������#������#�����@ �   �����V�?�����@ �   ;  ��a ����      	�    �    ���@ �   �?�X�      ��! �?�X  �`��@ �`���^��X��	B�����
�      	�    �    ��h  ��c�@ vj   �����  ?��� ch���'�D�'�H�'�L�'�P�'�T�'�X��T��X�?����\��`�'���'����D�  � �?������#�\����#�`'  ����#�d)  �� ��#�h�����������   +  ��`���`�    �    ����?������#�\3  ��`��#�`5  �����#�d������������   ������   �?����D����&� �&���P����"  �" ��H#  �`p�@ �`�#  �# ��L'  ��h�� ���$@ �$`'  ��ഀ���    �    +  �`p�@ �`�#�\�#�`-  ��h�� ���#�d�#�h��D�� ����P�� ��  ��`  �� �@ u�   �����  ?��� b؝��'�D�'�H�'�L�'�P�'�T�'��  �� �� �* @ u�   �'������� �    � 	     �� $@ u�   � @ u�   ��D��H/  ����� �������?����1  ��!� � 5  ���� � ��l   9  �� ��'�����;  �`��@ �`���L�?�����  � ��  � ���P�?����p����@ �`�"� �`�"��`�"��"���襠 ��#������#���������#�@��1      ��`�  � �$� � �$�� �$��$�� ����#�@��P      ����  � �&` � �&`� �&`�&`��p����  � �"� � �"�� �"��"���੠ ��#������#���������#�@��      ��`�  � �$� � �$�� �$��$�� ����#�@��#      ����  � �&` � �&`� �&`�&`��`����@ �`�"  �`�" �`�" �" ��p����� ���"` ���"`���"`�"`����#�@�߹      ����  � �%` � �%`� �%`�%`��p����� ���&� ���&����&��&��#�\��`����� ���#` ���#`���#`�#`� @���  ����  ��!�  �� �@  9   )  ��!����������?�ؘ�����������@ �   �� �    �    ���@ u   �  �    ��`����@ �`�"  �`�" �`�" �" �ܯ   ��T�&� �&���L����&� �&���P����"  �" ���@ t�   � �    � �����  ?��� b؝��'�D�'�H�'�L�'�P�'�T�'�X�'����H�* @ t�   �'����Ā� �    � 	     �� <@ t�   � @ t�   ��H�#`��D�� �    �      �!  ��`T��D@ t�   ��   ��`��\�@ �`�"  �`�" �`�" �" ��p��X�� ���"` ���"`���"`�"`����#�@���      ����  � �'` � �'`� �'`�'`� �'����Ģ �'�������H����    � 4   ��`����% �@ �`�"  �`�" �`�" �" ��p��X�� ���"` ���"`���"`�"`����#�@�ܠ      ����  � �#` � �#`� �#`�#`��� �'������'��������'�������H������   �    �'�������H��@�    � K   ��p���.���P�@�@ �`�"  �`�" �`�" �" ������+���Ĥ@�� ���"` ���"`���"`�"`����#�@��a      ��`�  � �"� � �"�� �"��"����* ��T��	�� ������#�@�ܬ      ���+ ��L���  � �$  � �$ � �$ �$ �����'�������H������   �    ��`��H�.`��ĸ��' �@ �`�"  �`�" �`�" �" ��p��\�� ���"` ���"`���"`�"`����#�@��_      ����  � �%` � �%`� �%`�%`���5  ���� � 9  ��! � � ��z   �'����D� ��H@ s�   �'��� �'����������@
�    � �   ��Ȓ����%   ��H���� �'���'�������H��@�    � j   ��������� �,���P� �@ �`�"  �`�" �`�" �" ������.���ĺ �@ �`�"` �`�"`�`�"`�"`����#�@���      ��p�  � �$  � �$ � �$ �$ � �������� ���"` ���"`���"`�"`����#�@�۬      ��`�  � �"� � �"�� �"��"���������- ��T���� ������#�@���      ��������.`��L���  � �'  � �' � �' �' �����'�������H�� ���   �    ������'��������������   �    ��Ȓ���ۣ   ��H������'�������H@ s.   �  ��D� �`�'���'�������쀦��    � j   ���������@	�*���P� �@ �`�"  �`�" �`�" �" ������- ��Į��� ���"` ���"`���"`�"`����#�@��:      ��p�  � �'` � �'`� �'`�'`� �������� ���"` ���"`���"`�"`����#�@��!      ��`�  � �"� � �"�� �"��"���������/ ��T���� ������#�@��j      ������ �+���L�@�  � �$� � �$�� �$��$���� �'�������쀦@���   �    ���@ r�   �����  ?��� c@���'�D7  ���(�?��;  �`��@ �`�?��;  ��`���  � ��  � ��	B  �`��@ �`��@�?�������虢�  ���0��	N�?��  ���� ����ء�	��?��  �� ��� �    �    �'���      ��a8����+���D�@�$� �$�������'�����+  ��`��� ���   �    � �   -  ������ �    � _   /  ���8�?�Ȱ �'���    3  ��`�����@�#�`��`��9  ��!@��	��������	\��ȅ��@�?������`�'�����  ��`��� 	���   �    �'��� 0   �����  ����� �����H��ؙ����?�����������P�#�`��`�#�`��`@ x     ��!8���@�#�d��d�#�d��d  �������#�h��h�#�h��h@ 	W   ��ȵ��@����*���D�@�#� �#����� �'�����%  ������@���   �    � J   '  ��਀����    � C   )  ��!H��D�%@ �%`-  ���H/  �����-���D�@�&� �&�� �'��� (   ����� 9  � ��  � ���D��ؑ�����ؑ�	��?�������Й�	N;  ��a8���  ��!P��	��#�`��`�#�`��`@ N   �����	�����* ��D��	�"� �"����� �'��  ��`��#`����� ���   �    #  ��`���`�    � <   �'��� 1   %  ���X����,���D���� �����X�#�`��`�#�`��`  ��`h  �� �@ q�   +  ��`���`�    �      �� �� @ q�   ������'������'���    ����'������`�'������'������'�����;  ��`��� ���   �    �����  ?��� ch���'�D�'�H�'�L�'�P�'�T��D�'����H� @ q|   �'������� 	�    � 	     �� p@ q\   �  �k   ��H� @ qg   �'��  ���`����� �����\�?����̘ �'��  ��a`����� �����@�?����̠ �'��#  ��ah����� �����D��葢F�?����̦��'��)  ��!h����@ �`��	J������L�?����̬��'��/  ���p����  � ���P��詥R�?����̲`�'��5  ���p����� ����	V��൦�X�?����̸ �'��;  ��ax����  � ���\��聠^�?����̒`�'��  ���x����� ����	B������D�?����̘ �'��  ��ap����� �����H��虣J�?����̠ �'��#  ��ap����� ����	N��।�P�?����̦��'��)  ��!h����@ �`���T��豦V�?����̬��'��/  ���h����  � ��	Z��ཧ�\�?����̲`�'��5  ���`��H�.���D�@�  � ���@��艡B�?��  ��a`��H�*���D� �`�`��	F������H�?��� �'��� �   !  ��!�����@ �`���L�?����̤��'��'  �������  � ���P�?����̪`�'��-  ���h����� �����T��ر�V�?����̰ �'��3  ��ah����� ����	Z��н��\�?����̶��'��9  ��!p����@ �`���@��؉�B�?����̐ �'��  ��ap����� ����	F��Е��H�?����̖��'��  ��!x����@ �`���L��ء�N�?����̞��'��!  ��!x����@ �`��	R��Э��T�?����̤��'��'  ���p����  � ���X��ع�Z�?����̪`�'��-  ���p����� ����	^��Ѕ��@�?����̰ �'��3  ��ah����� �����D��ؑ�F�?����̶��'��9  ��!h����@ �`��	J��Н��L�?����̐ �'�������襤�P�?�������୥�T�?������`�'������"���� ��e   �      ��a���L��P���X  ��ᐵ�����赦�^��T�$  �$ #  ��a���L��P���@%  ��������������F��T�$��$�� �    � �����  ?��� b���'�D�'�H�'�L�'�P�'�T�'��  �� �� �* @ o�   �'������� �    � 	     �� �@ o�   � @ o�   ���-  ����� � 1  ��!�� � ��|   ��D��H��L��P���5  ����� ����	��?��7  �����'�����9  � ��  � ��	R�?�����;  �`��@ �`��	V�?����p����  � �"� � �"�� �"��"���豠 ��#������#���������#�@��6      ��`�  � �$� � �$�� �$��$�� ����#�@��U      ����  � �&` � �&`� �&`�&`��p����  � �"� � �"�� �"��"���ൠ ��#������#���������#�@��	      ��`�  � �$� � �$�� �$��$�� ����#�@��(      ����  � �&` � �&`� �&`�&`��`����@ �`�"  �`�" �`�" �" ��p����� ���"` ���"`���"`�"`����#�@�پ      ����  � �%` � �%`� �%`�%`��`����� ���#  ���# ���# �# ��p����� ���#` ���#`���#`�#`� @���  ���  �� �@  "   )  ��!��������	��?�������������T���   �� �    �    ���@ o	   �  �    ���@ o   � �    � �����  ?��� c���'�D�'�H�'�L�'�P�'�T�'�X�'����H�* @ n�   �'����Ā� �    � 	     �� �@ n�   � @ n�   ��H�%���D�� �    �      �!  ��`���D@ n�   ��   ��`��X�@ �`�"  �`�" �`�" �" ��p��T�� ���"` ���"`���"`�"`����#�@���      ����  � �$� � �$�� �$��$�� �'�������H��@�    � 5   ��`����.���Ē@�"`�� ���"  ���" ���" �" ��p��T�� ���"` ���"`���"`�"`����#�@�ֿ      ����.`��ĸ��  � �'  � �' � �' �' ������'�������H�� ���   �    �'�������H����    � 0   ��`����- ��Į��� ���"� ���"����"��"�����/ ��P���� ����p�#�@���      ����+ ��L���  � �$  � �$ � �$ �$ ������'�������H������   �    ��`��H�.`��ĸ��' �@ �`�"  �`�" �`�" �" ��p��X�� ���"` ���"`���"`�"`����#�@�؛      ����  � �%` � �%`� �%`�%`���5  ����� � 9  ��!�� � �ն   �'����D� ��H@ n   �'�� �'�������쀢@
�    � f   ��Ȓ����a   ��H���� �'���'�������H��@�    � L   ��p����, ��Ħ��� ���"  ���" ���" �" �������  � �"` � �"`� �"`�"`����#�@��      ��`�  � �"� � �"�� �"��"����������- ��P���� ������#�@��O      ���������.`��L���  � �'  � �' � �' �' ������'�������H�� ���   �    ������'�������쀤����   �    ��Ȓ�����   ��H������'�������H@ m�   �  ��D� �`�'���'������������    � L   ��p����/`��Ė�	�� ���"  ���" ���" �" �������� ���"` ���"`���"`�"`����#�@�ՙ      ��`�  � �"� � �"�� �"��"�������� 	�*���P���� ������#�@���      ���������,`��L���  � �%  � �% � �% �% ������'��������������   �    ���@ m1   �����  ?��� b����'�D;  ��`���  � ��  � ��	F  ��a���	H�?�������𕢉L  ���������?��  ���� ��  �!��  � ��	R�?��  �`��@ �`���V�?�ؐ��!  ��!Ȓ � %  ����� � �ԧ   )  �� ��� �    �,   ��赠 ��?��+  ��a�-  ���ؽ����?�Ȯ �'��� !   ������@ l�   �#�h��h�� ����� ���艡	F��	B��Б�	D�?�������
������L��������R1  ��!੥	���ȭ��T�?������`�'�����7  ��਀�����   �    �����е����?��9  ��!��?��� �'��� �     �� �� � ����*`  ��ธ�
�  � ���  �`��@ �`�����?���������+�#  ��`��@�� ���"  ���" ���" �" ���1  �� �� �@ �`�"` �`�"`�`�"`�"`����#�@��      ��h�  � �'` � �'`� �'`�'`��Ȥ���� ���"� ���"����"��"������؍��H�#������#����ذ���#�@���      ����  � �&` � �&`� �&`�&`� ����#�@��      ��x�  � �"` � �"`� �"`�"`� �� �#�@��      ����  � �%` � �%`� �%`�%`�����𕢉L�#�h��h�#�h��h@ 
}   �;�p  ������
���#�x��x���#�|��|�#�|��|���@ ]   ���������T������p���V�?�����������X�?��5  ��������    �    ����#�\�#�`  �� �  ��`�������@ l   ���� �'�����  ������@
��M   �      ����� ��������\�?��  �� �� � �����B��D�#@ �#`  ��ഀ���    �      �� �  ��`�@ k�     ��พ��� ��  ��a   �� ����@ k�   ��D�� ��  ��aP  �� �@ k�   �    !  �� ��� �    �      �� �  ��al@ k�   �����  ?��� c����'�D�'�H�'�L�'�P�'�T�'�T� @ k�   �'������� �    � 	     ��!|@ k�   � @ k�   ����$������D��H�$� �$������L��P�%`�%`�����T�%�����    � �����  ?��� c����'�D� 
   ��D�`�'����D@ k�   ����'�D��D�� ���   �    �����  ?��� c����'�D�'�H��D�� �    �    ��H�    ��H�� �    �    ��D�    ��D�'���    ������'������ �� ���   �    �����H�#���D�    � �����  ��H  ��!��?������?�Ѐ� ����?���?���а���?��� ���� �  � �-��@�@ ���#��
��'@ ���@ +� ���'@ �@���@�����$� 
 � �����Ȩ �?�ж � �?�� � �'@�� $� � �����ȉ�B� ��?�Ѐ�@6� e��@!� ���$� a��@�����н����+�D������D0  �* �  �@�2 �
 �#�D��D            � � �@�  �& �-�� �& �����ॠ���ȩ� ���ȁ�D���T��	D���@��������#�h��h�#�h��h�;�H��H� %��@���F�  �-��� ��?�З� ?�����J�%����%������؝����@�& � �& ������������؍��P���B���B���P���Ʃ���#�x��x�#�x��x�;�H��H��@�� � {�?���+�D��D0  �`�/`�* �@�#�D� q��D   � ���2� 0�� ��Ѐ� 	�    �* 
� �� 
� � �  �� "� ��������Ё��^      #� b���� a�� >�� 	�    �* 
� �� 
� � �  �� "� ��������ȁ��\      3� M���� L�� >���� H��^2� &�@!  ��!���ȁ�
F      3� 	�����Ё�
F      #�   ����� 5���H�!��  �� 4� ��	T�� 5�?�Б�	X����?�������  �!��  � ��	@� �?���� � �'@	�# 	�%� ���� �  �#@	�&� �& �-�� �& ��������ȿ� !��  �����	^�?���@��@2� ���������@ Ř �?����Ё� >�� ?�����  ��x�?���?�������
@      #� 	�����聩
D      3� � ����Q��^�2 � �2   ��!���
N      #�   � @ �� �� !�A��  ���� ����
T�    � 8�@	�� 5�� 4��
X      #� &��`� � � � @ �� �� !�)��  �� $�&�� %�� $�#�� %  �  �" �a��@ �`�  � ����\  �� �� �� �!  �!��  � �������� �/`  w�aH� 	��      �� �� �� � �� 5�� 4��
J      � �� 2� +  �%  ����� �� �'  ����� ����� ｣�)  �!��a��@ �`�  � � 潤�T� � �
 	�� 	� � �  �� � `���� �
 	�� 	� � �  �� � J��`� T�/`  w�b4� 	��      �D �X �t ޔ-  ����� � ���/  ����� �� ���� ��� 9  �  ��" �a��@ �`� ���	^  �  �������� ��� ����^  �"�  � ��   �b�@ �� ��`� ��� %!  �  �� �!��  � �� ��� ����H#  �b �@ �� �%  ����� ���`� ���΀�`� �/`  w�cX� 	��      ޴ �� �� ����� �
 	�� 	� � �  �� � �� 2� -  �'  ����� �� �)  �!��  � ��� h����+  �a������ ���@ �`� _��Z����* �2 �;�H�����H�* �2 �;�H  �b�?���@ ��H�`�?���?��@ ���� @ ����' �� <$� ��`  ��b������@  ����� ����B� .�?��� ��?�6� ���  ���� &�?�������蕢���#�`��`�#�`@ ���`� �?��� &������   ���'���  ��������𽣈�!  �" �  � � ����������#  �b �@ �`� ������`� �/`  x�aL�@	��      �� �� �� ��� >�� ?�����  ��X�?�����#��?�ض � ��ܪ �@��@��� ���#  �b@�@ �`�� ���?��������@ A� ���?��#� �� 4�  ��؀� "� �  � �� � � � � �  ��@2� ��؀�@4� ��؀� "� �  � ��@� � � � �  ��@"� �������������^�6��* �2 �� �;�H��H�  � "�5`#� ��@&� %� � � ��@&� �� �?`�&�����$� �� �  ��4�>@
�.�
� 	���2� �� �  ���?@�.����2� �� ���  ���� 2� U�� ��@2� � !� �' �� 2� %� ����{���ހ� � 
�� 2�   ��t��ؐ"8�  �p� "�   �����k�� ��b8�@ �g�`��@
2�   �� �   ������8�� �����P      #� 	  �������@ 
�� �� !�Q��  �"@�  � �L�����J�����@2� � ����D���^��@2� �� �� "� �� �' �� "� 	�� ����;�H��H��@�� !�3��  2� =�� �� � 	%� �� "� ���� �� 2� 3�� ���� �?��  �b@�@ �`���ހ� � 	�?��������@ 
�� �� !���  �� 2����� �� 
2� ����� 2� ���  �"8�  � ��  �� !��	��?��������@ 
g� � ��?��2� �������   ��� ��'��2� ��耐 2� ���  �"8�  � �� $�� %��	��?��������@ 
M� � ��?��%������;�h��h@  ���l�� !��@� ��  � ��@&� ��������ؽ��H� 
��	Z�����警	V��0��ұ�	^���R��V���Z$ �?���� ��@	&� .����@	2�   ����� "� ����  �b@�@ �`@ �'�������@ 
� �� !� ���    �"8�  �?�艡Z� ��
�      � B�?��  �b@�@ �`@ ��'�������@ 
 � �� !� ���  �c��@!$3��@&� 0� #0$3��@2�   ����� "� ����  �b@�@ �`@ ޔ80������@ 	� �� !� z��    �"8�  �?�艡Z� ��
�      � �?��  �b@�@ �`@ Ɣ80������@ 	͘ �� !� b��  � �' 	��@$�   �  �� �� �"(  ��b0������D!  ��"8#  ����\�b@  ��h��F  ��`�� �#�x��x���#�p��p��� ?�/`�@��	L�@ �`  ᡤ��?�衦��  �bp�@ �`��	V�� ���"X���V�  � ��	Z���  �bP���Z���P�@ �`��	B  ���@�@�@ ��B�`��	H��蝣�H���N�? ��<��R�?����Z� �?�����@ o� � �?���� �/ � �%� �� � ���2� ������   ��	�'������� >�� ?�����  ��p  �  �!���#�"@��H� �� ���  � ��@�?�������� X�  #� �b��@6� T  ��𽧈���%� �'@��@2� ��^  �"8�  � �&� �&��  � �� /  ���  ᭤�֐"��  �   �b�  ����� �����  ��  �"��  �   �b��@ ���V���`��ܱ�	\��,��2��	Z�� ���L���Х��R��ę����� �����L��	P��̵��H��P���D��	T�@ �`��T��	D���D��	J���B��	X���\���V���R��ʽ�,���ڥ����&� � i�&�  ��@6� + �!  ����"x�  � ���T�?��?���� + �#  �@�c��@/� �@  �&� �@	?���@
�&@ �&`��������B�<`�$c�� ����#  �b�%  �!  �  �∠"�����  ���� �� ���#�`��`�?`'  �›`��	F�@ �`)  ������ ����0�"@�/`�@���^���\-  ���@�@���B���H��ֽ��D����� �����\���Z��	L���R���F���R��H���V��Z�  � ��
��H���\�@ �`��ܹ�ޭ��ܵ��V��Z��Ľ�&���̙����&� �&��� >�� ?�����  ��x� �* �2 � �;�H��H�?���?������ �
 	�� 	� � �  �� 2�   �� c��@�"@��
�      � ���@  ����  ��"H���@�"H���N      3� S�� >��	@���^��	�� M���^  ��"P��
�      9� ��  @ G���  ��bH��	�  ���\��X� :��	@!  ��"��  �� !� ��
�      +� +  �@ 3���#  ��bX� ,��	^  ��"`�bp�@ �`��	J'  ���x�� ����	J���-  ���h�� ����́���      '� �;�h��� 	� � 
� � � 	� @ '��  ��h@ ��l�?�����#�@ ��  ��  �� !�� >�� ?�����  �㿀� � �
 	�� 	� � �?��  �� 2� ������� d���^�. �2 �;�H  ���H�"��  � ����      9�   ��;�h��h@  W��l  ��b���@  ������	����   �
���L��	N�#�h��h�#�h��h�* � 
�;�H� (��H�☁���      9�  ���!  �  ��"��"��  � ���T  ��b��@ �`���T���ځ����#�h��h�#�h@ ���h�?��������   �
��* � 
�;�H��H�?�����@ ��#�� �;�h��h�;�`�
 	�� 	� � �  ��`�� 2� �� >��� 	� � 
� � � 	� @ ���  �� >�� ?�����  ��@�?������ �;�h��h�;�`�
 	�� 	� � �  ��`�� 2� �;�h���^      �   ��"�����      =�   ��O���^�M�b���h�2 �� "� �/  �  ���Ё���      =� F/  �  ���؁���      =� 
���^  ��#@�  � ���H�?���3�� >  �c��@ �`��	N  ��!  ��� ����N�#��  ��	@� #  �c��@ ��	F�`  �#��  ���F���Z� '  ᵦ�Z��  ���	J�b����P�b����@���й�	@������ �����څ��D��ą��ʅ��Л� !��  ���F���F��F��H�����\�������      =� G%  �5  ���0�� �����@  ��#8�  � ��D  �#�  ၠ޹��^  �c������D�� ����	J�  � �@ ��	@�`  ���� ��@��  ቧ	D���J�#��  � ��	N  �c��  ���D��D� !  ��"荧�F����#  ���Z���ʍ��J���ڝ����@ �`���ʝ��Ɲ��X���N��	@��N��X���\���H�b�����^�������      =� 	)  ���l@ ���h'  ��������^�# ���^�?��-  �+  ��bȬ�H�� ������^������      9� F#  �5  �������      9� 
���^7  ���@�� �������?������ >9  �#��  � ��	H  �#�  ��  � ��H�c��@ ��	L�`  ����� ��	@��  �#��  ��@���Z�   ᵦ�Z�#�  ���	D�b����J�b����L��ʹ�	L�����  � ��ڝ��P���Н��ĝ��ʏ� -�� ,���@���@���@��B�P���\�c����      9� �)  �%  ���0�� ������  ��#8�  � ����+  ��c ���܁���      � 7���ҽ�	\/  ���� �����J5  ����� ����J7  ���� ���@��9  �#��  ���F�   ����� ���F��	@��  ၠ@�c��@ ���J�`-  ���艧	D������ �����B��ȱ�X��	H���ȕ��؉�ʉ�	Ɲ�N��Z��	D���\� 6���Z��	\  ���� �����J  �  �#��c��@ �`���D�  � ���J  ���� ���N����D  �#��  ���H� #  �c���	N���N'  ���	@��ر��X��ā�	D�����葠��@ �`��đ�	���Z��	H���H�  � ���H���Z���\���N� ̽��^�#(����      9� �/  �  ��"��;�����+  ��cX   �@ �`���^�
��* � 
�;�H��H���@-  ���0/  ���R�� ���#�������8�#��������� �����@5  �������F������@��ځ��� D���!  �#��  � �  9  �#��;��@ ��;�`�� !������^��  �  �   ፧	F�#��  � ���F  �c��@ ��	J�`  ����� ��	B���  � ���B���J  �#�  ᱠؘ#��  ��	F���J�  � � ���@������`�  ���� ���Z��	D���č��ځ�Ɓ�	¹�	L��H���@��@��H� A���\���^  ���� ����	B#  �!  �#��c��@ �`��	L�  � ���B%  ����� ��	F����L  �#��  ��	@� )  �#��  ���F���F� �;�p���H���!  �#��  � ��̹�	B�  ���Z��	L��ځ���  � ��́�	ȁ�N���@���@��N@ P�?��������p��X�  � ��^� �#�p��p�#�p��p@ B��  ��P�� ������      � 	�;�h��h@ *��l5  ����� ��^��h��l@ "��  �� >�� ?�����  ��h9  �#��  �?��������Z� ;  �c��@ ��	B�`  �#��  ���B� ��	L  �c��@ �`��	F���L  ����� ����	B  ���?�𽦉F���F��𕦉N���޽��^���̹�	N���ޕ��L������ �����̅��ʅ��P���B��Z��P�����  �㿀7   �?��!  �#�. � ������6� 0 � ���6� ��	@� ���6� ��	@� `� ���B� ���� 	��	B� ���F� ��F��	F� ���F� ��	F� ���F� 0���F� (��F���F�  ��F���F� ��F���F� ��F���F� ��F���@��	F� ~��F���� M�� ���� H �  ��	���	@� 0���F� (��F���F�  ��F���F� ��F���F� ��F���F� ��F���F�  ��F� X��	F� )��Ā��� � �  ��	���	@� H���F� @��F���F� 8��F���F�  ��F� X��	F� ��Ā��� � �  ��	�� X� ���� X���� 	�� ��&���@	�    ���� 6���� P�� &� 2���� 0����   ����� �  �?�������	B�� &� �������� �  ��F  ��#`��	ƶ' 
�6�  ��bh�����	@"� 	� 8� H���H� @���H���H� 8��H���H�  ���H� ��	H�@�� &� ��́�L� ��J��ʁ����  ��@!   �. %�H�����@� � � �  @ �  �����  !� ��@� ����?�����������@ n   �
 �, ���%  ��,�Ā   @ �������   @ >�����灠 �@ ������だ �@ 6������   ��P�?��!  � ����5   �. � ���� � ��.���@� �   �� � �   � �� ����� r)� � �  ���&� 	�  4� E�� � ��@8� A�� �  ���4� �� �    � $����    � � (���� 0���� � � (��B� 0��J�?��� ���	@� p���D� h���D���D� `���D���D� X���D� 8���D� P���D���D��Ā�� � 	   ��	D��Ν��΁���� @� r������	D���ĝ��Ν���� @���ȁ��΀��"� h��@� H� e���@4� �  � ���&� � �� 	�� 4� � � ��@(� � ��� � V� � T� ��	B� H�� 4� ��F��Ɖ�D���'��� ����H�������� ����J�>�� ��ʀ��� )� � ���B���� � @� 5��D� H��	F��F��	F� /��F�  �  ��	@�/ � Љ��D� ȉ��D#  �ah���D%  ��h���� 8�������	H'  ��h��	�������@��Ā� � ��|&� 	�`6�/`�'�����@�'��� 
���/`�'�����@�'������ ����@�����  � � � @ O� ���   +  ��@���   �@�/�����+3� �� � 	   �"�@�'������'����������偠@   �* 
�;�H�����H   �* �
����;�H�����H�㿀�?��!  � ��  ���#���c��� %�B4� )��B#� �� � �#  �� � [#   �. ��@� 	�� � � (��	D�?��?��� P���� � � � @ 	� � �   #?� �� 6� �����  � � � � @ �� � �   �� &� � #��� � d#� �� � 1   � ���@�� �* #� �� 2� �  �& ��@"� v�  ��	D� ���D� ���ȑ��H� n��ȑ��D����	���c��& �"@�����	H6� 	� `� p���J� h���J���J� `��J���J� X���J���J��ʕ�	J� T���'  � �4��"#��@#?� �. #� � �'��� #?��������  �?���������'�荠B�4���	������  �! ���F��� P��	J� H��J��	J� @���J��	J�  ��J���J� 8��	N���N� ��N� 0��	J� $���J  ?��� �
�	�  �?������������B�& ��	Ƒ2 �*   ��ap  ���p���F� P��	J� H��J��	J� @���J��	J�  ��J���J�@��J�����J�����  ��@!   �. %�H�����@� � � �  @  {�  �����  !� ��@� ����?�����������@ �   �
 �, ���%  �����Ā   @  f������   @  ������   @  ^�����だ �@  �����߁� ���@�?��+   �. ���!  �"`%� ��@� %� ��@6� ��	@��@� E�  %� ��@&� 	�  � 0���J� (��J���J�  ���J���J� ��J�?�𕠉J�  � 2��J  �@���
@�'���'��� ���" 	�2`�� ���� ����?������� 6� ��D��ą�	@  ���p� @���J� 8��J  ���ȕ��J� ���N� ��N  ��" ���N�  ���N��	��	N��	J� 	���N������	��ʁ�J�����  ��@�?��+   �. ���!  �"�%�@��@� %� ��@6� ��	@� N��@%� ��@&� 	�  � 0���J� (��J���J�  ���J���J� ��J�?�𕠉J�����	J"� :��J���J� 6��J  �@���
@�'���'��� ���" 	�2`�� ���� ����?������� 6� ��D��ą�	@  ��� � @���J� 8��J  ���x���J� ���N� ��N  ��!p���N�  ���N��	��	N��	J� 	���N���J��	��J�� 6� ��J�� ���ʁ����  ��p!  �#p�?��� �� � ��  � ��@� �� �    � �����  �>`�'����`� ����� ���B� �   � � ?  ��@���     � ����    �. ���� ��� � �   � �����	B�?��������   � ��	B� x   �� � z���� u   �/�����?� �*�  ���'���'��������� ��	B�6 � �"@� 8�2 �
`���	�� �" �'���'��������J���D� (��Ɖ��F  ��	D�?�����"��'����葢	F� (���ȉ��H�������� !�'�ؗ3 <  �+ 
  � 
�  �  �'���?�����  �" 	�'����艡�J���         �����?�����  �" �'����蒂`�B  �?��� 0�  �?���/�܉�	D��ܐ� �    ��
B      � 	   ���         ��@�    �� $�� %�?������ ����������C  �'���'������ �����聠B      ��؁����  ��������@������?� �
 
���
� �* 
�� 	�    ���@���� � 	� @  �   ���   ��@   !  � Т. �H�!���@�>� 4� �&� &� �&��!��@8� �&� �&��&�� ��   ��!|��@� � �� � 0����H�����@
"� � H� 8��ƅ��� ����Ɖ��� P��ʅ��� �����NH�!���@4� L� �� � ��	B� ���D��B�4`��� 0��	J�'������ 8��	L�����&� �� �2��
���"@
���� 1���#� � H�� *�� +��	P��Й�ʙ��� P��	N����� $���̡�	P����� P��	N�����&� �� �2��
���"@
���1� ���D� � X�� *�� +��	P��Н�ʙ���� `��	D���� 
���̡�	P����� `��	N� ���̙�	L���̡������� >��̀�@� �4`�� ����>� �>�� =�  �"��*��$@	�&� �� ��@�  ������ ��	F�?����J�����ā�	F�?�聨
V      � 
   � ��
V      �    � � �?�� �'� � �   ��c8@ 	�   �� � � �  �� ��   �@���&� � 
�&��� � � �� ��� ��  �>� �>������  ��P  �!�?�и' @ ]y�?���������?�耧 (�/ �c�?��  ��c� 	��      � d   � d  � ` 4  � � � ,   � � | P �  d !P "� #� $� %� &� ( (� )x * *� +L +� ,� -8 -� .� / /�!  �  �cp�"��'�� � � �'��@ <� %  ��?�����'  ���`�?������ +  � !��%bH@ 	!����� 2�/  �-  ���`�� 2�   �  ��a�� @ ]!�   � !��""H  ����  ��x�'��  �� �"��'��� � � @ �?��  ���`�?�؀��� #  � !���$bH@ ������ 2��/  �%  ���`�� 2� )  �  ��a�� @ \�� )  � !���%"H����?��  �〔 �'��  ��"��'���?������"�   �
��* � 
�;�H��H��
D      � ���� ������  ��c0�@    �
��* �`� 
�;�H��H  ��b��?��  ���`�?������ #  � !���$bH@ ������ 2��/  �%  ���`�� 2� )  �  ��a�� @ \�� )  � !���%"H  ��c-  ����@ �'�� �'���`�?��  ��c`�� 	2�   �  ����� �?��� x�  � �'���'��  ��#`�� �   � "�~�#�H@ ������ 2�z/  �#  � "�u�$bH)  �'  ���"��'�� � � � @ |�'��-  ���`�?�؀� 2�   �/  ����� �?���`x�@ �`�?��  ��c`��`�   � "�T�"�H@ W����� 2�P/  �  � "�K�#bH%  �!  �#�����'�� � � � �'��@ Q)  ��#`�?�؀� 2� /  �+  ��b�� �?����x�� ���?��/  ���`����   � "�*�"bH@ -����� 2�&/  �  � "�!�"�H!  �  �c��"��'�� � � �'��@ (� %  �����?��'  ���`�?������ +  � "�
�%bH@ ����� 2�/  �/  � "��%�H  �c�  �����'�� � 
� �'��@ �    ��#`�?�؀� 2�   �  ��b�� �?����x�� �� ����?��!  ��#`�� � %  � !���$�H@ ����� 2��/  �'  ���`�� 2� +  �  ��aԔ @ [� +  � !���%bH  ��"�/  ���'�� � 	� �'��@ Ӑ   ���`�?�؀� 
2�   �  ����� �?��� x�  �� �� �?��  ��c`��`� !  � !���$"H@ ������ 2��/  �#  ��c`�� 2� '  �  ��a� @ [�� '  � !���$�H-  �+  �c�����'�� � � �'��@ ��    ��#`�?�؀� 2�   �  ��b�� �?����x�� �� ����?��  ���`����   � !�u�#bH@ x����� 2�q/  �  ���`�� 2� #  �  ��a�� @ [x� #  � !�b�$bH)  �'  ���"��'�� � � � @ i�'��-  ���`�?�؀� 2�   �/  ����� �?��� x�  �� �� �?��  ��c`��`�   � !�@�"�H@ C����� 2�</  �  ��#`�� 2�   �  ��b� @ [C�   � !�-�#�H%  �#  �c�����'�� � � �  @ 4�'��)  ��#`�?�؀� 2� -  �+  ��b�� �?����x�� �� ����?��/  ���`����   � !��"bH@ ����� 2�/  �  ���`�� 
2�   �  ��b$� @ [�   � !���#"H!  �  ���"��'�� � � � @ ��'��%  ���`�?�؀� 2� )  �'  ����� �?��� x�  �� �� �?��+  ��c`��`� /  � !���%�H@ ِ���� 2��/  �  ��#`�� 2�   �  ��b8� @ Zِ   � !���"�H!  �  �#��"��'�� � � � @ ��'��%  ���`�?�؀� 2� +  �'  ����� �?���`x�@ �`�?��+  ��c`��`� /  � "���%�H@ ������ 2��/  �  � "���"bH  �  � ����"��'��� � �  @ ��'��  ���`�?�؀� 2� %  �!  ��"�� �?����x�� ���'���'��%  ���`���� )  � !�w�%"H@ z����� 2�s/  �+  ��c`�� 2� /  �  ��bL� @ Zz� /  � !�d�%�H  �c�  �����'�� � 
� �'��@ k�    ��#`�?�؀� 2�   �  ��b�� �?����x�� �� ����?��!  ��#`�� � %  � "�B�$�H@ E����� 2�>/  �'  ���`�� 2� +  �  ��b`� @ ZE� +  � !�/�%bH  ��"�/  ����'�� � 	� �'��@ 6�   ���`�?�؀� 
2�   �  ����� �?��� x�  �� �� �?��  ��c`��`� !  � !��$"H@ ����� 2�	/  �#  ��c`�� 2� '  �  ��bt� @ Z� '  � !���$�H-  �+  �c�����'�� � � �'��@ �    ��#`�?�؀� 2�   �  ��b�� �?����x�� �� ����?��  ���`����   � "���#bH@ ې���� 2��/  �  ���`�� 2� #  �  ��b�� @ Yې #  � !���$bH)  �'  ����"��'�� � � � @ ��'��-  ���`�?�؀� 2�   �/  ����� �?��� x�  �� �� �?��  ��c`��`�   � !���"�H@ ������ 2��/  �  ��#`�� 2�   �  ��b�� @ Y��   � !���#�H%  ����#  ��?���c�'  �� ����'��)  ��#`�'�䀐 � �?��+  ��b��}�?��@ ������ 2�y/  �  ��b�� @ Y�� /  � !�o�%�H  �c�  �����'�� � 
�'��� @ v� ����?�ؑ2 �� "� !  �@ 	������ȁ�
B      #� !  �  ��"����F�;�`�#�p��p�#�p@ 	���p��@��`���@      3� !  ����   ���'��!  ��#`�� 2� )  �#  ��b���Ё�
�      =� '  �%  �� �� ����=� �?���"���Ё�
�      =� -  �+  �`x�@ � �`��x�� �� ����� 7�?��/  ���`����   � "��"bH@ ����� 2�/  �  � "��"�H  �c�  �� �'���������'��2 �� � �?��@ 	������ȁ�
\      #� ���!  ��"���	B�;�`�#�p��p�#�p@ 	}��p��@��`���@      3� ������#   ���'�����-  ���`�?������   � "���""H@ ܐ���� 2��/  �  � "���"�H#  ��c  �#��@ � �'���`'����Ȧ���'���+� ��������и  � �?���  � -� ���&� �� �>��'c���`$� �� �  �`4�>��.���@2� �� � ��2� �� �  �`�>��.���@2� �� ���  � �� � �� 2�   ����   �@�'��  ���`�� 
2�   �  ����� �?��� x�  �� �� �?��  ��c`��`� !  � !�}�$"H@ ������ 2�y/  �#  ��c`�� 2� '  �  ��b̔ @ X�� '  � !�j�$�H-  �+  �c�����'�� � � �'��@ q�   ��#`�?�؀� 2� ���  ��b�� �?���?��  ��#`�� �   � !�L�#�H@ O����� 2�H/  �!  ��#`�� 2� %  �  ��b�  @ XO� %  � !�9�$�H���  ��c�@    �
��* �`� 
�;�H)  �#�� ��H�'��+  ��c`�'�䀐 � �?��-  ������Ё���      =�   �/  �� �� �#��=� �?��  ��b���Ё���      =�   �  ��x�� � ����x�� �� ����� 9�?��  ��#`�� �   � "���#�H@ ������ 2��/  �#  � "���$bH)  �'  ����"��'�� � � � @ ��'��-  ���`�?�؀� 2� ���/  ����� �?���?��  ���`����   � !���#"H@ ֐���� 2��/  �  ��c`�� 2� !  �  ��c� @ W֐ !  � !���$"H� ���%  ��'���   �* 
�� 	� �'��� �  � �� 
2� �� 
� � 6� �* 
� � �� 	2�   � � �� 
"� � � �� 2� 	)  �)  ��#�  � �'��� �'���"Д � @ �� �?��-  ���`�� 2� ������� �?���?��  ��#`�� �   � !���#�H@ ������ 2�|/  �!  ��#`�� 2� %  �  ��c � @ W�� %  � !�m�$�H� ���)  ��'��    �* 
�� 	� �'��� �  � �� 
2� �� 
� � 6� �* 
� � �� 	2�   � � �� 
"� � � �� 2� 	-  �-  ����� ���'��� �'����Д � @ Q� �?��  ��c�@ �`�?��  ��c`��`�   � !�1�"�H@ 4����� 2�-/  �  ��#`�� 2�   �  ��c8� @ W4�   � !��#�H%  �#  �`����'�� � � �'��+  �@ $� �c�@ �?���`�?��+  ��c`��`� /  � !��%�H@ ����� 2�/  �  ��#`�� 2�   �  ��cT� @ W�   � !���"�H!  �  �  �"��'�� � � �'��'  �@ �� ���� �?�����?��'  ���`���� +  � !���%bH@ ܐ���� 2��/  �-  ���`�� 2�   �  ��cl� @ Vܐ   � !���""H  ��(� ����'��� �'�� @ ΐ  �?�����%  ���`�?������ )  � !���%"H@ ������ 2��/  �+  ��c`�� 2� /  �  ��c�� @ V�� /  � !���%�H  �`0��А �'�� 
� �'��@ ��   ��"���Ё���      � �?��  �`x�@ � �`  ��x�� �� ����� !!  ��#`�?���� � %  � "�x�$�H@ {����� 2�t/  �)  � "�o�%"H���-  ��8�'�� � 
� �'��@ w�   ��?�������`�?������ #  � "�Z�$bH@ ]����� 2�V/  �'  � "�Q�$�H-  ����+  ��?���`@� �'������'���?��  ���`����   � "�?�#"H@ B����� 2�;/  �  ��c`�� 2� !  ���� @ VC�   ��c�� @ V>� !  � "�(�$"H'  ����%  ��?����D� -  ��'����`����'�䀥�� �?��  � "��""H@ ����� 2�/  �  ��c`�� 	2�   ���� @ V�   ��c�� @ V�   � "� ��"�H  ����  ��?���`H� %  ��'����`����'�䀤�� �?��)  � "� ��%"H@ ����� 2� �/  �+  ��c`�� 2� /  ���� @ U�   ��c�� @ U� /  � "� ��%�H  ����  ��?���`L� ����'��  ���`�'�䀣�� �?��#  � "� ��$bH@ ǐ���� 2� �/  �%  ���`�� 2� )  ���� @ UȐ   ��cȐ @ UÔ )  � "� ��%"H  ��"�-  ��?����P� �"��'��  ��c`�'�䀢`� �?��  � "� ��"�H@ ������ 2� �/  �  ��#`�� 2�   ���� @ U��   ��cؐ @ U��   � "� ��#�H  ��"�#  ��?���`T� �"��'��)  ��#`�'�䀥 � �?��� r� "@ w����� � p/  ���`�� 2�   ���� @ Uy�   ��c� @ Ut�   � "� ^�"bH  �  � ��X�"��'��� � � @  e�'��  ���`�?�؀� 2� %  �!  ��"�� �?����x�� ���'���'��%  ���`���� )  � "� <�%"H@ ?����� 2� 8/  �� 3� "  �  � `����'�� � 
� �'��@  <�    ��#`�?�؀� 2� #  �  ��b�� �?���`x�@ �`�?��#  ��c`��`� '  � !� �$�H@ ����� 2� /  �)  ��#`�� 2� � !  ��c�� @ U� � !-  ��%�H/  ���`���� 
  ��#`�� �   ��c`��`2� �������� >�� ?�����  �㿐� �+�D��D�  �* �'�H�@�2 �'�L�� �#�H� ��H�+�D��D� �`�*`�* �@�#�H��H0  �+�D��D�  �* �@�2 �#�D��D�� "� �� �+�D��D0  � �*`�* �@�#�D��D�� � ±.   ��a�� 	��      1� 2h 3( 3���`2�  �  �+�D��D�  �*#��@
�#�D��D�2 �
 � �
 �+�D�* ��D��H�*#��@�#�D  ��c�@    �
��* �`� 
�;�H��H� ���D� �;�H��H�?����H���   �
��* � 
�;�H� ���H��`2� !��H�� 2� ��H�+�D��D�  �*#��@
�#�D��D�2 �
 � �
 �+�D�* ��D��H�*#��@�#�D  ��#   �
��* � 
�;�H��H� i��D  ��#(�     �
��* � � 
�;�H��H�  � � [���V��`2� #��H�� 2�  ��H�+�D��D�  �*#��@
�#�D��D�2 �
 � 	�
 �+�D�* ��D��H�*#��@�#�D  ��c�@    �
��* �`� 
�;�H��H� 7��D  ��# �     �
��* � � 
�;�H��H�  � � )���X��`2�    ��+�D��D�  �*#��@
�#�D��D�2 �
 � �
 �+�D�* ��D��H�*#��@�#�D  ��c�@    �
��* �`� 
�;�H��H� ��D�#�  �� :� �� ;���ځ� >�� ?�����  ����   ��  ����'�T�/ � 
�'�D  �!ؐ&��'�H� �&�@ S��'�X�� � �'���'��������� �*`�*`�@
�&�	�'��� �" �  �" �.��  �� 6� ��X  ���� � ���@�� ��X�@�� �#@ �����`����#`�� ��D� A�    �� @�� &� �  � � 	�� <�� � .�� =�  �"���`���.�� � ��X� �  � ���� ��	F��X�&���
�� ���H��������	J�`��`���&���콧�L�� 6� �/ ��X���� ������ ��	N���&��`��󽧈P�/ ����@
�"@ � �� ����"`  �  �  ��`H�?����P� X�?�� � ?��c�����'�� ����  ��'��� @�?���� � � �'��� � �  ����'�Ā� 2� �  � �  ���'������ �'��� �'��� � �  �'���,`������� ���,`�  � �$`�"0�  � ��	\  �b(�@ ��@�`��h��������^�@�'`��ƴ&���\�#�x��x�" �@ �`��^���� 6���  �����;�x��x�;�p��|@ ��;�`�����	R�;�h�  �#�x��x�#�x@ ��x�����	V��h��������`��V�� �#�p��p�#�p��p��� ���ޞ�d�,`����d������� �;��+��" ��d�"� �@���� � �:@����� "� ����,`��d��� �>`����      7� � �� $� N  䀐 �  �  � � ��h�.����� 2� ����� "� �� @ �  ��	��h� � �#��  ����h�"������&����h����� 2� ���� ��`�,`��d�@
�@ ����@� �"@ ��d���� ����
�
� �#� �� ����� "����,`��`2�   �  �" �  � ���ހ� "�   �� �  ����;�`@ 0�;�p��p������`  �b�@ �`���J      #� �  ��$`���� #�  �&���@� �.���h���&���h� �@
�@�&���h� 	�&��&���h���&�����@�@���&����&� 	�� ��h� �&��@����&��� 2� ]  ��% �.�� � �&���h� �� "����`����`������X�@�' �*��.��/ ��X����@����
� =�&��� ���� ;�%� �%���Ā� 	"� .� �  �"���`���.�� � ��X� �  � ���� ���P��X�&���
�� ���R���������T�`��`���&���콧�V�� 6� � ��X���� ������ ��	X���&��`��󽧈\���&@ ��� �&`�`�� &��Ľ� :��Ţ@�`@���@      � ����$`�"�� �'���$`�"��'���,`��h� �� "������� 4  ��;�h��h��l@ ��  
�� !  �"(��  �  � ����      '� ��^�� #  �b0�@ �� "�`��	^�,`��h�`�,`��D��h�����H��H���ʝ�^�#�p��p�# ����#�h����h�'��� �" 	�,`��h�#�h��h�"�  �b �@ �`@ U����� !  ��0�� ��  ���,`�,`� � ������������T�&��'`�&����Z�"� �"��� 6�����h  ��`@� $� �$@�  �  �� =�"��  �" � �-��@���  � �@ �`��	X���`��� ���@�� 6� �$@�� &������$@�*`��Ȗ�	�"� �%��"��� 6��ݽ� <��T�� � đ*   ��b|� 	��      >� >� >� ?�  ��`@�,`� � � �  � ���D�&��&��� 6�����Ȁ� 2� �� �  �"0�"  ��H�" �"� � ��"�  ��`@�,`� � � �  � ���J�&��&��� 6�����Ȁ� 2� �� ��� >� �� ?�� ?��H�#��#� ��`�"� �"����� ���ޘ �# �# ���� ������� ���R�������T�������,������� 6� 	�� ���� ���V��������� 2� �� ���H�"��"��� � a��� � ��И �?��?��?��?���@�#?�޶&���\�#?��#?��#?� 4���.��$`�'`�,`�� 6� ���  �� @�,`� � �@����������H�&��'`�"�ޝ�\�"��"�����"����� �����R�&��&����6�����Ȁ� 2� �� �����#���H�#�   ��#@ ��0�#`�����H�"��"���H�#��#��� � ����ȩ� ��#��� ?��H�#� �"�   �"0�"���Э� ���H�"��"���H�# �# � �    �"0�"  � �" �����  � �
����
2� �  ?� �* �� 	2� �  � ���   � ���"� �  ���"� �  � ���   � ���2� �     �* ���	"� �  � ���      �* ��@
2� �  � ���   �;�H� �� � ��H  ��`�� ��	B   � �#�H��H���� 
�:�� �"�5�� 
�:�2� �"�����#����   �㿀!  �"`#   %� �� 2� ����?���. �- �� � 4����  ��	B����� H   �&�6�?������ � �6�2� �6��?���. �- �� � !���+  �� �    � ��@���� �/ �    4� ��'���?�� *� 6�/ �. � �?��� ���� 	��	B&� �. �    � �?����������  �/�����+1  �� � 
   �. +� �@�?������ ���	B�!)�'������  � � �?���������/�����+1  �� � 
   �. +  �@�?������ ��ہ�	B� ��'������  � �?������������2 �㿀!  �"�#   �. )� ���&� �  �?������  ��B�    �'���'�������B��ª ��
D         �    � 0����'������- �@�'����������  �㿀!  �"�#   �. )� ���&� �  �?������  ��B� $   �'���'�������B��ª ��
D         �    ���� � 0���H         -� 	���� ���H         ;� ��D�'������- �@�'����������  �㿀�/�����2 �* �6 �+ � 	  �b��@�> ���c�� �� 
8� � 
� ��@:� 	� � @  )� ��@�'��� ����'������� �����  �㿀     �� &� 0x w��#�?� �?��� 8� � 
� ��@	:� 	� � ���� ��@�'��� ���� �'������� �����  �㿀!  �#8�?��)   �. ���+� ���� �� �  ��B�    6� �  � ��B��
B         �    �� 6� �  � � (������  �㿠�����  �㿠�����          ?�              T�I�%��}@      ?Tz�G�{?�������@               ?�              ?�              ?�      ?�              ?�              ?�              @$      <�      <�      ?6��C-@              ?�                      ?�              @!�TD-?�      �       ?�                              ?�      ?�                      ?�      ?�      =�|��׽�        ?�      ?�                              ?�      ?�              ?�      ?�              ?�je
\\?�      ?�      @               ��      A.��    @D�     @k      @;      @q      @T�     @      @�@             ?�      ?�              ?�      ?�              @      ��      @       ?�              ?�      @      �      ?�              ?�      ��      @P      ?�      ?�      ?�,�>w�a?�Y���t?��Eu��?�Xl��?���2�Ѣ?��[Q?�B���-�?�r�<}Q{?�[�o�u?�ԇ1h��?�;�b��?�8znub8?�kEe�|�?����?�҅��?��
1�?�<�d�?�q�7:��?��4��?�ަL4"?�
!�.*?�N`a�-?􆢵�<�?����6*'?���v�,�?�4+V�O�?�oG6�'�?���HT)?��o�!H?�$~�:U�?�b8�U"%?���f;�?�߲<e/?�u��_t?�_�VBg�?��s��?���6�Nb?�%��L�?�hٛD��?���B*��?��w6?�77����?�}���NP?�đ���?�f{]�e?�U�>%]?��kUy��?�蟙Zӭ?�3��O�?�v��^G?���K��?��݅R�?�g�.W�K?�� ��i?�-J�|?�X����?����2�?���3{�_?�P.�?�?�������?���aZ'?�Pv[nE@?�������        �q��S[]<�s�u�e<a��K���<��.J�a
<@:'�{S���9D�:��/���6����A�׊v<�[L{Ih�<�n �d<<��u�J��<��~��s<��3�@��<�语U<�GT�A�<��j�1��<�'!�6Y���:�B��u�6�a��<��	𞼼^�i0�x<H�z��<s����b�<}C���B⼔�	�YW㼀z��<�<��,��<�2LFG�<���0��^����~@�����	�Y4���4�dV�k�:h<����nG��z���$YW1mӼ�w��/<p]�y~��L�2�<�����<���V�K'<����l�g_ǁ�~���[|��<||F�q򾼓YI]�3��/nۍA�<�����1<���4]́�b�^0���uXO~T�;<�=�z-��<�e�PH�<��M�H<�<u���Iۼ��7Cyz�<���[7<�# im�2����OK\<�����̏���#�(�<��􆤶�<���-ء�<�HS�        ?��P    ?��    ?��    ?���    ?�M�    ?��8    ?��/    ?�c�    ?��    ?��B    ?�r�    ?��X    ?���    ?�*�    ?�v�    ?��    ?�B    ?�L+    ?Ɏ�    ?��^    ?��    ?�I�    ?΄    ?ϼ    ?�y
    ?�    ?Ѭ    ?�D    ?��    ?�q$    ?�F    ?Ԛx    ?�-�    ?��    ?�Q�    ?��!    ?�q�    ?� �    ?؎�    ?��    ?٨    ?�3v    ?ھ    ?�G�    ?���    ?�Y/    ?��    ?�gS    ?��?    ?�rj    ?���    ?�z�    ?��y    ?�?�    ?���    ?��    ?�    ?�@�    ?�(    ?�1    ?���    ?�<A    ?�zL    ?�    ?��h    ?�2|    ?�o?    ?㫳    ?���    ?�#�    ?�_:    ?�x    ?��j    ?�    ?�Jn    ?儂    ?�M    ?���    ?�1    ?�j     ?梯    ?��    ?�>    ?�K    ?炽    ?�    ?��2    ?�(	    ?�^�    ?��    ?��    ?� �    ?�6    ?�k�    ?��    ?���    ?�
~    ?�>�    ?�s    ?�    ?���    ?�A    ?�A�    ?�t�    ?�i    ?��    ?�m    ?�>�    ?�p�    ?�X    ?���    ?�?    ?�6c    ?�gS    ?�    ?�ș    ?���    ?�)    ?�Y    ?��    ?�U    ?��    ?��    ?�E�    ?�t�    ?�N    ?�Ѿ            >6��
/��>@�ZE1M�>Z�f�]�)>Mc�a�M�>W!Ukޟ>c�S�Vy�>k��8[ �>oY"bϙ�>[��֫��>P+j��>1����>q�O<r��>r�okԋ>|O�C�>>0~�'>\��C��>z��O�8>z�v_�E>-��|�:>V�vI���>y�)��N>c�[�=->|��I��>>w MDu>�v-�c>�Zan�a.>�R>
Q�>�a��0H�>���U��o>�ԙ��2&>m��$��z>r�F⿒K>����o��>l��C��>���tܤO>������>�O�g|��>xŇ��>|�,�i-�>�#���W>l���]�>D���:��>~_��8i>��T��>�<�h�>��+j���>�GK�+�>�]A���>��Fɉ�c>�<�A�4>|�8�G�>z2����L>�P�W9�>�r�/�r�>�O��Kh>�T�J�>�*yOc�>�T<�sµ>��R�I�>n���>�a�$�H,>�����>F/��<>��޴<� >�z�Ʌ	�>��')��>�m�,H�>�T,ٙV>{ϸ5qT>���Y��>�@�� >��F⿒K>����|>���)>���q�6>sLN����>Yj(iU�~>���5�c>��	K>���y��>��A�A3>���Rv_|>�b��|��>����xܯ>�����y>�&�\�=W>p�g��g>���[{�>�Od��>������>}���ٴE>f ��C�>�h*˧2>�U�����>�v	�Ү>��l̫>�I�%��&>�q��2>�����>���o��>��9Z*�>s^d5��w>zT�E�]>��[Iin>�s�,��>l�~m��>�tضj>�\4
�m1>��<8��>��&bƿ�>�Q �Ho>�I�%��&>�O�:�/>�]A���>�Y�0�>�g�����>pCW�%��>w ��U>~Dg+�>�lMNUD4>�Qa�l>�l�T[p>�;n�d2>�y�ʩɫ>�����7>aw�3b��>�ʾP��?�-V�?�      @6      ?�      @�      ?�.B��9�?�.B��  =�9�5y<v@�.B��9�?�      ?�      @�@     @�      ?�.B��  =�9�5y<v@�.B��9�        ��      ��.B��9�g�FFԗ��.B��9�?�      ��      �D      �n���Y?�.B��9�<g�FFԗ?�?;�s?�\���s�@Q�     ?�.B��  =�9�5y<v�������       @�.B��9�?�Ge+��?�պ��/n?�����?����7&?�ܽ����?�����bl?�Ї��O?�Ɂ>�j?��ԉ�3�?ǹ{K�[?Ȱn⇜(?ɦ��l�&?ʜ#@2y?ː�R�`�?̄��t.n?�w�� W6?�j���M?�[u�,��?Нŗ�cb?ы���x?�x7 W�F?�bw7��?�J�6¯
?�0��Q�J?��	��?��A���?��`Kc��?زM9J%?ٌ�EMk?�d���#�?�:��\l?���N��?��SC,P?ݬga�O?�@�T?�e~��0�?�%]��ҩ?������?╎Y0�1?�E��7�?��?����?䗏�&��?�8�{�?�Չ��?�mf9#��?� ��xF4?�k�]1^?�з�M?���W��?�!�TD-?�%��%?�O8d��?��p�C��?�|W�o�?�nW�O
�?�$�D�U�?���|�A�?�sҁ��?�.4�?�Ng'z�?��GS�?�ӏ,[��?�� 9�?�K���?�_@0�?���D?�b���6?�p�U�:%?���A�m�?�myjM�?�O��	?�jl�3S?���P��G?��kz�`?�-pA��?�[T�sQ�?�L��?���e��?��x���?����g&?���D�?�6����?�oo3��?��PRN`?���ڽ?��s%HW?�Ʃ+�?�AMD	L|?�`�,sj?�}�c���?��!:�PS?����0�p?�ǌ~ޱ�?���{�e�?���C_�?��@1�?�^� ��?�$���j!�L�v�v�mq���<|���d�<X�V4<f;�(<a�#��X�PT�,=<{Z�b�<SG�����<ws�g��<L��4�<`��ʅ<!{��嫼Y[���&<ld�4Y~<hf� )�e<h�n<���<v.G9�e<c�t���pw��m���ic�D�rؼu��<U���bVd��@��zrWq <��*���t<v��\+$�<{m�t��<y�Ɉ�
w<��	�W� <zᇱ�P@�|��p�L4<����*<z+"/e�j9��8*#�}[I_cI�R�����5�Y(�(zf��p�s����<�7�<~ϋI&D�<rA���X���t��R<`�K��ʼv�o�軺�x�M%���<����7@�{�b)ӹ��[�^z<��&3\�h��a�����i6�3�z+V7,�<���:ъk��c�Ej�n<�z��3ؼRb�;]��<p�z�˽<�4=����<gT��>�<�i��� ¼���#�p��+/�^U �r�p�?��YR?
�ӵ<�Fj���<��v(ևH��f��_��<�+-X���<�%L�;��<�y��aռ�,w�\<��;5�tm�DA��?�<������<y�.�ļeg��Y2Ѽ��>�'�U�l�zc�A�<�4����6��W���oG����}�����;<x��ȝ�<������]��Q�;Qʼ���α���_`�\s��z�j�3*����.�����9Q�㼗ѫ���<�#�� �⼒��Dy(缉W���|��"���W��*<����Hh��ށbF��Ť����D��s��b[�K�Y�$�U�Ű���E��O��
=u��+'^)����zWͨ�lM2&u��IJ�$�i�&��D��*@� 㷵cH�� �����$� ��?;�s� c�	�� &�|;e���WU� 2��b�������sXB���~pbdl��*�����e�����NApˏ!���S�mc���+Ͽ���-��?6�����Tt��v��b��ל�P��ț�GpԿ�t&��3��!f���^���I�F忿������,��2�+�ng���+d����������Q4�?6���u2~Y���x��Έ��{t�Aڿ�6��T�����O�7����M�It��n�X\�P��.B��9���8��Y#��5�x��ڿ��5�K�:��K҈����ۘ��;K��n\��Gu����[���D櫿�7�Nr*���k�Pl��t
PA���s"?��ӏ$7}��_�KE���I�Y��b������
@,-���'&ο�rP�������>N�h��73XN����I\���*�����t&��3���'�j�ÿ�T�ʥc ��ȥ*�Iſ�>��0�緍�D5#��2Xט�3��E��Ա��.B��9��2.&�xW��=���#ſ�P(������ib4ے���@�<���v��T��߳X�zH����'&ο���ETɿ��)RH�п�s�CV�����;��֊�>�j��"�8�ؿ��Rw31���ib4ے����'�|�ϙl��y��7�e^{�ʓ�<����#�eQ�¿ſ@kT=���e�������'�|���'c�F���3^]YI����] ~�������:������C��A]��DD�� VX�XG        ?���x3 ?�
0�b�?��Ҋ�kL?�'n*��?R��#?��0p���?�RZ��V�?̏�ǚ�"?Ϲm^>+?�g\���?����1?�a��^�?�ѽ�X	�?�9����?ؚ3��B[?��#쿘L?�D�{̏c?܏�ǚ�"?��j�ġ?��_��?�%R����?�r�%*�?�T�����?��_^p@�?�y^��?��3O�?���V*?���Fr�?��]�>�?�*-&[ū?�@L5�-?�.B��9�?�*W�m��?��
�P?�]PV�Y?��#쿘L?�ӗ�78?�$�?�٦7O�?�R@���x?��Q�z?���T��?\jȈ?�/�p4�?����Sj?��},�?�=�a-m�?��z�?��_^p@�?�;qcÀ?�< �� ?���Wh޳?�)��Pw?�vZ�9?���h���?�Q.�=`?�SЈ���?��$�W?���(2?�%�s�VO?�i��U<U?��8���?������?�.B��9�?��Mk4�?�&����?��P'���?��u��?���]�8�?��),j?�X�R���?��A��3?�%f��?��)�#s?��{���;?�F��Q�?���n�<b?�����-�?�T�ઊ�?���* ?�����]�?�R@���x?��]�*�?�������?�@�Q�"o?��|q�1?�ؤ�t��?�"r�2ZW?�j�?}?��.���N?��3h�N�@ �y���@ @_��,�@ a��b@ �q����@ ��?;�s@ �uX��@�;��@Z8Ӓ��@��z�@�n���@�FF$�@7��
��@k���U@�C��V@ϝԱ 5@�Ζ��@.�7L@\��&��@��>%t@���ӿ@��Ӟ}@Q.�=`@4�8.��@]?��@�+1�Q@���@�N�D�@��3���@�׻�@A	���@d�o�@��t5�@�9MH@��V��"@�=�Ҝ�@RI?@.B��9�@mH5*U@�k��z@�ɓQeJ@{:k��@W�.|9A@�6�,@�h��Z@�B{s�@)ԅ��@[.�o��@�_VV]�@�tw=��@�z��;(@	}�ѳ�@	A�o�b;<�7eN��<��>�1E;��־񫼍�w��\�<�<�����<�wx;.`<�:^}�<�uH99K����{Ƽ���)�)�<��	삖N<�{��[�<������⼭;�)"Q\��vҒ�d�<r�\fѼ��V5����>�+�9<����w���vw��"��ěk�5���G��x���ל�&��[m(�Zj<�S��wμ���y	c���Ӫ/�<��U�=0R��y}���м�	;�� n��~��V�༁f
H�8�<�;�U�������y���K*{�4<���ޱ�<�(Q�����9逻C/��:c��0<RF��z�Z<���S\I���nĳ�!<��vϧX<R����;<� ��kԼ��~�vB���>}��iм��AW������;9�?��"�C�ƼCj�W<I&����<���ŏ�<���֟0<��O�x�<�S�f�;��־�<|1lW�<��}_�PN�l�_�|�<�rh��s�<����Z_�<�oէ��<��"jtC���ěk�4�rI����<��Ȥ߸�V��5.�A�aD7\r�<��|&9�<�釳�w�<N][X.��v��y���ގk�&"���:�&�<h乨o�J6�ƃ���2�iO�1���t����3��wX�z��;9�?�y��J�aM<xOHQ�<�`eQ\���ݝ�*����V��������N�g��Y$�Y<z�Ȥ߸�b#��eJ�y�lE�>�<h�(σ�<RJ�;w�Zd��tx<h�鳊iy<r�'�
�Ƽ~�ݝ�+<`�:_Ƒ�ofPf����f)$$q��k����r<a#,��<!��L��W���D�<P�:_Ƒ�T�qs0<Tx�W̷�Wi�,xB̼a�~�g�:��v`�=�L�u6"�2|���        <3>?��#<H_2\[�ͼYّ����6x b<cw@}��[���on<m�LN.&�d���C@�l��d��<,�>��7�x�͹^��<B����<t#c���x�l�K�r�9߻���J��!\�|�D�E�x�t���C@�pFvVظ��s(��8ü|��Q@� ��Y�3 ���3hv<~�,����d���F��<o����fڼ���g�H:<�/0�<1=�=7a��a�7P�M
�CYUh?q�<z��;9�?<{��+��1������4�����Z��!\<P�g%f�z<s�|zdd<��b$�K����S`t�s���?�&<{��0��������<�����'�<�p ߋ <�}LTO<�	��cѼ�%o�ʫ�<��,����<WQ� �����Ϝ)��6 l@�B�?R�`p��c�+�Y�<��A+ռ��M<s#w<px��4x��Z&\��<����;󼉈���'�<{�}��[<q����Y�<xQs�1�<���;9�?<�V�3a�<�!H����p�y��-漚��c�漘A���0(��^�׼��N�r�7<��}ޔX��7��:��g�e/r<�!�E�����]�2��1��?м��:G%B�}�iH�|<�o�hI����iM����S`t�<�L����<��X��９�#��b༛Ν����<d���|_%<��R[<���2����<�U1�l�<d��M�<����L"<�ѣ�H��<�����?��<{��;m<��V5�<�-7�?s�<J��������+j��%o�ʫ뼨�-8h���u!�Sd�� ?�����H�IN��<��A����<�GC)�0�<��!�	�X�������t�9N��<�ۛq��n��L������@�[ז���M<s#w�������<���Zy�G�#u�(<���5�^<��G�8^�����"<����T<�|~�"M>��\�X�ּ����<CAș5�J<�Rn�_��<��o�M֎��F��km�<���;9�?<�	�7MG����h1�꼫i��e�<�2$-��<��f�`��<����ܤ<�7S�q�<��~���ط�d��t&U��K<�?�fp�`���U���<�⻎P<r+�����xZ� ?�4
|�(?�)p�p?��@7M?}��6?�L.��?��Wo�2?�|���$?�vS*w��?�pkߞ�?�je$\��?�d>��*�?�]�t�5	?�W���g�?�QM���?�Jl�:y?�C��<��?�<�ó�n?�5�he��?�.��S��?�'f���?� 0�d�?��)i>�?��	Ň;?�	/�8\~?�T�}�?��A0/&?�����?�ϧD��?�!Ov�?� a��O?ç̓?�)��?�s>�=@?�_T�6��?�J�K*D�?�6��֥?� �I���?�
�Z��?���>��^?���P�(�?�Ʒ�Y?�k���?��/q��?�~N��{J?�e?>@@?�K����?�1���|?�Pr}��?��l�R��?������?��J���.?���}?�[���?�o9 ��;?�Q���^?�3��݁?�([}P?���1��?���X�?�U:AN?��Ab��?�̵&���?��Cs�-?�=}R��?��h�/�?駵�je?�Zg���?��xM��?�Z]� ?�i�w��?��1�m]?���	�O?�i��U!?�o�vx?渘���]<�[k;tb<�-F��;�g�?M:�L�>(�e$̘��e�3+�z!r�(�x�[�u@��|¶a�>����6ܴ<���$<v�
��(�����(<n:>�Լ��g�$70<�=��W��y��B�b:Ҋ4�<�ͤ?��<��!_VՂ�b�/����<{���K��en�L�<��rv,�<GPV:��<�<���������r�K�#��ñ�Um
J�Aм�/��T><b��>�e���&K�<�<�9z��X���B�5F�<���/ȼ����.�h3�rw��R7�V`���ck<_��w漎-�~g6ļn���+��<T�dwm�5<�$�+^\�<������c�p5+피�b6CK�7<�4�w��a<~`�0���<��+���<���P�*<��9�1�<d�+�:��dj�H^4b<z�ѡY#��A����B�a��;��������������(<s�Ȍ�<TZ<Ǐ��<X�yGz<q�V���<��j�ֶ�<i�8^ǒ����졖i��� �y<�"�̟��������,�p��
�;�<�c�>�t�<s8���ݼm��(޼ls��*�h�h'�όh�<�%����<qZǆ���?��1,]f�?�i�����?���M��{?�f'�ƉY?��Oϡ&�?�ba�-��?��]�ZML?�^B�*�S?��/��?�Y��<�]?��c.��D?�T�W}"?��R���?�O�$�_?���)ze?�I�a%��?���N�a�?�C�u��?���X���?�=Rz�8?͹�_���?�6R��H�?β���?�.�����?Ϫ���w?�Q\�e\?�� ��d6?�Ha����?��}dƸv?�>R�6?Ҹ��>��?�3���?ӭ�i��?�&���?Ԡ�= ?��h�z?Ց�����?�
)�u?ւ�8��?����:U?�qUvB?����mN?�^z�iI?�Ԥ�t�/?�Jk��F�?ٿ��?�4���?ک[c��w?��2?ۑ>0۬C?���@�?�wg�ў?����ԥ?�[�4va?��L2��?�>V�X*i?ޮ�tK�?ߎ��j��?�6)9ƙU?��?��Ķ�;?�|�_.�?��426WL?�P��x��?��B?� T�H�O?�YtV(+?��%�l�:?�N���8k?��F��a?���{5?�q��mY�?�����?�,��!�y?戊NK/<d}fkfˑ<%w'y�L<YI�*�r��lbo�5��f�C?��<Ts#��3���,\���<bQ۾=�<E�P�<��<[���S*�b�b˹S<j��4�<Y�=��}<h��a�U�Y�;W���<6��Ɇ��<i��j{�����f&�hhЛ�|k�V�Y�G�4�c. ��o¼2@�?9c��`��W,�f-�·�a]�P�2��y���Ǽy�
�ⴼk聵��<t`v����t��3N�<aU8���<~��0,< =U���<�{T}0<x#�k���<{5qU���<g�K�?��<[���3�}��DJ�<t+�N���f��1K�μ{c�ڿZ�<x��_��<tJ�vc&�v��>h?X<p�9� ���Z1;P�ͼf)>�<��z�B˙��~8�/l?�<a��u~���^�M=X&�b����<r�D�_<p���q���P������W��<�}<Y�P�- �����x9{���C�9�<�������<c^W.$�<r*?��Z<~��$W�μ��q�!j�<�kB	Z[�q��;��[�p�W����ljU< �s�Ŝ����aĈ0<\�;M��<�l�p�W���ݘU�$����vD��?�              G����   ��      �����   ?�      �����        ��������      �������       @	!�TD- ��� nND )� 'W� �4� ��b ��< C�A �Qc �޻ �a� $n: BM� �I .�	 ђ �� �) �>� �5� .�D �� p&� _~A 9�� 9�S 9�� �_� ��( ;� ��� � �/ �Z
 mm 6~� '�	 �OF ?f� _�- u'� ��� �{= 9� �R� �k� _� �] V0 F�{ k�� ϼ  ��6 �� �a^ � e�� _� h@� �؀ Ms' 1 V� s�� `�{ ��k        ?�      @       ?�      NFS=%d
 AMPL=%.15E+i*%.15E abs(AMPL)=%.15E arg(AMPL)=%.15E FREQ=%.15E
  error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 Nbre de termes cherches trop grand  %6d  %-+20.15E %-+20.15E
   TEST/ECART = %g   ON CONTINUE
  TEST = %g ECART = %g 
  FREQUENCE   FR = %g  TROP PROCHE  DE  %g
   DANS ZTPOW, N = %d
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 error : malloc failed!
 KTABS2= %d  FREFO2= %g
 IFRMIN=%d IFRMAX=%d IFR=%d FR=%g RTAB=%g INDX=%d KTABS2=%d
 error : malloc failed!
 CORRECTION DE  IFR = %d AMPLITUDE  = %g  %+-20.15E %+-20.15E %+-20.15E %+-20.15E %+-20.15E
 error : malloc failed!
 error : malloc failed!
 ZDIV= %g+i%g DIV=%g
     %g %g %g %g %g
    g_NAFVariable.T0= %g, g_NAFVariable.XH=%g, g_NAFVariable.KTABS=%d
  F1=%g ,F2=%g
   T1= %g , T2= %g, T= %g
 FR1= %g ,FR2= %g ,XT= %g 
  DIV= %g
    error : malloc failed!
 error : malloc failed!
 DANS ZTDER, N = %d
  AMELIORATION PAR LES SECANTES
 SEC: A=%g, B=%g, abs(B-A)=%g 
  SEC: F(A)=%g, F(B)=%g
  ECHEC DE LA METHODE DES SECANTES
    DIVISION PAR PRESQUEZERO
   ON CONTINUE AVEC LA VALEUR TROUVEE
    ECHEC DE LA METHODE DES SECANTES
    BEAUCOUP TROP D ITERATIONS
     ON CONTINUE AVEC LA VALEUR INITIALE
   POSITION SECANTES %g TROUVEE A %g    SANS GARANTIE
  AVEC GARANTIE
 
 %19.9E %12.8E
     ROUTINE DE RECHERCHE DU MAXIMUM :
  ERREUR FATALE
   PAS D''ENCADREMENT TROUVE
     OSCILLATION DE L''ENCADREMENT ?
   %12.8E %12.8E %25.16E %25.16E %25.16E %25.16E
  %12.8E %12.8E %25.16E %25.16E %25.16E INF
   PLATEAU DE LA FONCTION
    COURBE TROP PLATE
  SORTIE AU SOMMET DE LA PARABOLE
    CORRECTION MINUSCULE
   %12.8E %12.8E %12.8E
    POSITION TROUVEE A %g PRES
     TROUVEE SOUS UN PLATEAU DE LA FONCTION
    
%10.6E %19.9E %19.9E %19.9E
   error : malloc failed!
 error : malloc failed!
 DANS ZTPOW, N = %d
 %20.3E
 naf_zradyd - N N'EST PAS UN MULTIPLE DE 6
  error : malloc failed!
 error : malloc failed!
 DANS ZTPOW, N = %d
 OMEGA=%g, DELTA=%g ,COR=%g
 CORRECTION DE LA 1ERE FREQUENCE
    FREQ. DE DEPART=%20.15E, CORRECTION=%20.15E
    FREQUENCE CORRIGEE:%20.15E
 PAS DE CALCUL
  error : malloc failed!
 acos: DOMAIN error
 asin: DOMAIN error
 atan2: DOMAIN error
    y0: DOMAIN error
   y0: DOMAIN error
   y1: DOMAIN error
   y1: DOMAIN error
   yn: DOMAIN error
   yn: DOMAIN error
   lgamma: SING error
 log: SING error
    log: DOMAIN error
  log10: SING error
  log10: DOMAIN error
    pow(0,0): DOMAIN error
 pow(0,neg): DOMAIN error
   neg**non-integral: DOMAIN error
    sqrt: DOMAIN error
 fmod:  DOMAIN error
    remainder: DOMAIN error
    acosh: DOMAIN error
    atanh: DOMAIN error
    atanh: SING error
  : TLOSS error
  : TLOSS error
  : TLOSS error
  : TLOSS error
  : TLOSS error
  : TLOSS error
  gamma: SING error
   ��                                                  00���     <0���     H0���     T0���     `0���     l0���     x0���     �0���     �0���     �0���     �0���     �0���     �0���           �    GH    GTo��� �o���        �       
  �                 o���       �      �          8          �   	                   @	!�TD-        @(#)hypot.c 1.17 92/03/23 SMI   �             @(#)atan2.c 1.13 92/03/23 SMI   5��zJԸ?�!�TD-?�!�TD-@	!�TD-<��&3\        @(#)pow.c 1.26 92/03/23 SMI             ?�      @       ?�.B��9�?ο����!?�k�z�?���TG��?U؁�Vw�C@      @G`   >d��c��@Ge+��?��	�9KS?�wrB��@G`   >d��]߇@Ge+��?��	�:�?�wlP��?�av���?ԇP�&CA@(#)_TBL_exp2.c 1.5 91/05/22 SMI    @(#)_TBL_log2.c 1.4 91/05/22 SMI    @(#)cosh.c 1.10 92/03/23 SMI    @(#)sinh.c 1.11 92/03/23 SMI    @(#)expm1.c 1.12 92/03/23 SMI   ?�         5    ?�p��<��?S�E&�?�q�8$��?P?�ˌ��?�      ?�      @(#)atan.S 1.17 92/01/13 SMI    ?�      ��UUUUT�?ə���_*��I$�ʹ,?�q�rm���A��?n?����=���UUUU;]?ə��#G���G`Y��?�!�TD-<��&3\G��CWi@(#)cos.S 1.8 92/01/13 SMI      @(#)exp.S 1.20 92/02/15 SMI     @�.B��9�@�I�-0Q?�?;�s?�.B��9�?�.B��9�?�.B��  =�9�5y<v@       ?�      ?�      ?�UUUUU>�f�l���?Vj�%�,���A��k�>f7ir���?�Ge+��<�              F)>Y9���?�.B��9�?�.B��  =�9�5y<v@GGe+��>�      >0      ?�UUUU)�f�fJ7 �?�      ?�Y���t?�Xl��?��[Q?�r�<}Q{?�ԇ1h��?�8znub8?����?��
1�?�q�7:��?�ަL4"?�N`a�-?����6*'?�4+V�O�?���HT)?�$~�:U�?���f;�?�u��_t?��s��?�%��L�?���B*��?�77����?�đ���?�U�>%]?�蟙Zӭ?�v��^G?��݅R�?�� ��i?�X����?���3{�_?�������?�Pv[nE@        <�s�u�e<��.J�a
���9D�:���A�׊v<�n �d<<��~��s<�语U<��j�1�伖:�B��<��	�<H�z��<}C���B⼀z��<�<�2LFG�����~@�����4�dV��nG��z���w��/��L�2�<���V�K'�g_ǁ�~�<||F�q򾼝/nۍA�<���4]́�uXO~T�;<�e�PH�<u���I�<���[7����OK\���#�(�<���-ء�@       @ Y���t@ �Xl��@�[Q@r�<}Q{@ԇ1h��@8znub8@�����@�
1�@q�7:��@ަL4"@N`a�-@���6*'@4+V�O�@��HT)@$~�:U�@��f;�@u��_t@�s��@%��L�@��B*��@	77����@	đ���@
U�>%]@
蟙Zӭ@v��^G@�݅R�@� ��i@X����@��3{�_@������@Pv[nE@@(#)fabs.S 1.14 92/01/13 SMI    @(#)log.S 1.23 92/01/13 SMI             ?�UUUUUU?�      ?�      @       C0      ?�.B��  =�9�5y<v?�UUUUq�?ٙ���:?�J�?Ei�?�UUUUT�?ٙ���:�?�I#O��?��Z��c        ?���x3 ?�
0�b�?��Ҋ�kL?�'n*��?R��#?��0p���?�RZ��V�?̏�ǚ�"?Ϲm^>+?�g\���?����1?�a��^�?�ѽ�X	�?�9����?ؚ3��B[?��#쿘L?�D�{̏c?܏�ǚ�"?��j�ġ?��_��?�%R����?�r�%*�?�T�����?��_^p@�?�y^��?��3O�?���V*?���Fr�?��]�>�?�*-&[ū?�@L5�-@(#)sin.S 1.9 92/01/13 SMI      @(#)__cos.S 1.9 92/01/13 SMI    ?�      ��UUUQ�(?�b�̝��������?�UUUO[5�V�k�U%i>��9�)9@������c(?�UQ_z�@(#)__sin.S 1.9 92/01/13 SMI    ?�      ��UUUQ�(?�b�̝��UUUUT�?���*�u�K�>�㦗'�������c(?�UQ_z�@(#)_TBL_cos.c 1.4 91/05/22 SMI @(#)_TBL_sin.c 1.5 91/05/22 SMI @(#)sqrt.S 1.19 92/01/13 SMI    <`      CP      >@      ?�      ?�      ?�      ?�������     .�  Mg  k  ��  ��  �z  �f  �J 	 � 5R I� \� n4 ~_ � � �E �� �� � ��  �� �� �~ � �� �= �f k� h> y� �M �� �� �E �a ɉ �m �{ �� � � �� �T �� �* �5 � �, �N �� �� n. R 3J Q  �Q  �  �  Y$  �@(#)__rem_pio2.S 1.9 92/01/13 SMI               ?�      Ap      ?�_0m�ȃ?�!�TD-?�!�TD-?�!�T@  =дabc1=д`    =дa`  ;��.ps;��.   9{��% I�@(#)_SVID_error.c 1.35 92/03/25 SMI @(#)matherr.c 1.6 92/03/09 SMI  @(#)_TBL_ipio2.c 1.4 91/05/22 SMI   @(#)__rem_pio2m.c 1.9 92/03/23 SMI                  ?�!�@   >tD-    <�F��   ;x�Q`   9���   8z% @   6�"�   5i�            ?�      Ap      >p      @(#)ieee_func.S 1.23 92/01/13 SMI       CP      <�      �             @(#)rndint.S 1.10 92/01/13 SMI  C0      �0      ?�      ��              �       ?�      A�����  A�      A����� A�      ��    ��      ��      ��     @(#)rint.S 1.15 92/01/13 SMI    C0      �0      ?�      ��              �       ?�      acos    asin    atan2   hypot   cosh    exp exp y0  y0  y1  y1  yn  yn  lgamma  lgamma  log log log10   log10   pow pow pow pow pow sinh    sqrt    fmod    remainder   acosh   atanh   atanh   scalb   scalb   j0  y0  j1  y1  jn  yn  gamma   gamma                               ��      �            �                                 �                      8           �           GH      	     GT      
     G`           x`           �           �           ��           ��           �p           �h                                                                                            �           7 �L         	         ��            ��            ��   #         ��   -         ��   7 ��   P     A �x  	0     K I  T     U �$  �     ` ��  �     k j|   �     v t�  �     � ��        � ��  L     � k0  	�     � �  �     � �  d     � F�       � ]�  �     � ��        � �h        � �p        � Ȩ  8     � ��  `     � ĸ  �     � �x   L     i�   �     ��                ��  $ ��       + ��       4 ��       <         ��  D ��       K �       Q �        T ��       Y ��       ^ ��       c         ��  i �       p �x       v �<  L    } ��       � ��       � ��       � ��       � �@       � �8       � ��       � ��       � ��       � �P       � ��       � ��       � �X       � ��       � ��       � �`       � ��       � �h       � �H       � �p       �         ��  � ��   !    �         ��  � �   !    �         ��  � �(       � Vp        Vx        V�        Vh                ��   �H       & V�       - V�       4 V�       <         ��  D WH       J W@       P �h       W W8       ^ W0       e ��   �    l WP       t WX       | ��        ��       � ��       � ��       �         ��  � ��         � ��         �����      ��  �   P      ��  �   X      ��  �   `      ��  �����      ��  �          ��  � �h         �   8      ��  �         ��  � ��         �   @      ��  � ��         �         ��  �   H      ��  � ��         �         ��  �          ��  �   (      ��  �   0      ��  �         ��  �         ��  � ��         � �,                  ��   �            �      ��     �      ��  $ ��         - �         2   �      ��  7 |         <          ��  B   (      ��  H   0      ��  N �h         P����      ��  R����      ��  T   �      ��  ^ �h         f          ��  q         ��  |   x      ��  �   �      ��  � \         �   H      ��  �����      ��  �         ��  �   @      ��  �   �      ��  �   �      ��  �   �      ��  �   �      ��  �   �      ��  �   P      ��  �  �         � �h         �   �      ��  �   X      ��  �   `      ��  �  �         �         ��  �   h      ��  �   8      ��  �   p      ��  �         ��  �         ��  � ��          h                      0      ��     8      ��   �         %         ��  /   (      ��  5 �         = �          A         ��  F         ��  J          ��  O �         Z �         b   @      ��  e   X      ��  h   H      ��  k   `      ��  n   P      ��  q   h      ��  t   p      ��  w          ��  { �         �          �         ��  �         ��  � P         � �         �         ��  � �`         �          ��  �         ��  �         ��  �   8      ��  �   @      ��  � ,         �         ��  �          ��  �   (      ��  �   0      ��  �         ��  � ��         �          ��           ��           ��  	   8      ��     @      ��   �                  ��  !          ��  $   (      ��  '   0      ��  *         ��  5 �        <         ��  G �0        N         ��  U d         a �p         j����      ��  l����      ��  n p         r 	         v         ��  | �         �         ��  �����      ��  �          ��  �         ��  �          ��  �����      ��  �����      ��  �����      ��  � �         �   (      ��  �   0      ��  � �         �   8      ��  � \         �         ��  � x         � ��            0      ��     H      ��     X      ��   �         !         ��  ' �         .         ��  3   `      ��  ;   P      ��  C   8      ��  K          ��  P         ��  X   (      ��  ]          ��  b �         k   @      ��  t �         }         ��  � w        � w(       � �8   $    � w0       � w       � 0�  �    � w       �         ��  � �\       �         ��  � �|   "    �         ��  � ��   #    � �(       � �          �        �0        ��        ��   @             ��  ) �`         2         ��  7 C<         E C�         S����      ��  U����      ��  W          ��  ] C�         m         ��  t         ��  y D         �         ��  �         ��  � ��         � E�         �����      ��  � ��         �          ��  �   (      ��  �         ��  �         ��  �����      ��  �   0      ��  �          ��  � D�         �         ��  �         ��  � �8         ����      ��            ��  
   (      ��           ��           ��  ����      ��      0      ��  $          ��  ) G@         5         ��  < 4�       F �      M A�   (    X ��   �    ^ �  "    m �   t    t h�   �     FL   x"    � '�   d    � ��  �    � mp  X    � 4�   "    � 9p   �    � �x       � ��       � �L        � .�   d    � �p         � R@       	    "    	 �D  	�    	 =�   �    	# o�  X    	/ �  @!    	4 ��   �    	B 4�   l    	N 8�   �    	Z �        	p լ   �    	� (   d    	� A�   ("    	� E�   �"    	� w8      	� D�   �    	� B8   h"    	� A�   4"    	� �@         	� �L         	� #@   H    	� 1�  �    	� .�      	� $   �    
     "    
 E�  @    
 Dd   �"    
 *�  �    
(        
3 �|         
: F�   �"    
? 8$   �    
L >  4    
^ �l  �"    
b ��  �    
q &<   �    
~         
� ,�  �    
� ��  �    
� GH     	  
� �p  �"    
� �l  �    
� D�   �"    
� �   "    
� ��         
� �      
� 6<   �    
� ��         
� A�   0"    
� 'P   d    
� D\   "    
� ��  �     c�  0     @�  4     �D  	�"      �  "    % 3�   �    1 �x  `"    = ]p       I 6�   �    V ��        _ \8  �    j @D   `    } �d         � �  @    � #�   D    � D\       � #�   D    � �  �    � ep       � W`      � :8  H    � 0�   �    � r   X    � ��  �"    � %l   �     FL   x     J@        �X         % �h   X    = B    "    D B        M �l  �"    Q ��   !    Y �H       _ tx  X    k H        w B�  �"    ~ �l  �    � B�  �    � ��         � Zh      � ��         � E�   �    � 4�  �    � �f        � �        � 4�   �    � B8   h    � A�   4    � L@        ��   �     �        # G`       0 4(   d    = ��         D Dd   �    K ��  �"    P (|  T    ] F�   �    d 5�   �    p H  �    u ��       x &�   h    � ��         � N\  �    � �p  �    � �       � D�   �    � 4  x    � N@       � GT     
  � %   d    �     �"    � �x  `    � $�   d    � A�   0     �  X     ��          7|   �     �  �"    $     �    * ��   �"   example crti.s crt1.s values-Xt.c example.c modnaff.c naf_funcp naf_ztder naf_ztpow naf_ztpow2 naf_prosca naf_modtab naf_gramsc naf_zardyd naf_profre naf_modfre naf_frefin naf_proder naf_fretes naf_fftmax TWIN BF AF naf_ztpow2a naf_maxiqua naf_proscaa naf_func naf_maxx naf_secantes hypot.c sccsid twon1022 two1022 atan2.c sccsid PI_lo PI tiny PIo2 PIo4 pow.c sccsid two53 log2_x B0_hi B0_lo A1_hi A1_lo one zero B0 A1 B1 E1 A2 B2 E2 A3 B3 E3 B4 E4 two E5 _TBL_exp2.c sccsid _TBL_log2.c sccsid cosh.c sccsid ln2hix ln2lox lnovftx ln2x sinh.c sccsid ln2hix ln2lox lnovftx expm1.c fminx fmaxx sccsid ln2lox ln2hix exp__E lnovftx invln2x q1 p1 q2 p2 atan.S constant exit x pio2hi pio2lo big tmp one N0 q1 p1 N1 q2 N2 p2 q3 N3 p3 p4 p5 p6 _TBL_atan.c cos.S cos_return casebase exp.S xflow ln2_32hi ln2_32lo constant TNaN huge exit ln2_2 ln2hi ln2lo S k x invln2_32 S_trail threshold1 threshold2 invln2 ln2_64 subnormal half tmp ln2 one zero twom54 twom28 twom18 t1 p1 T1 S2 t2 p2 p3 primary ln2_onehalf p4 two p5 fabs.S log.S constant small exit ln2hi ln2lo log_0 one_third two52 large_n TBL half one zero quick_cran log_neg A1 B1 A2 B2 A3 B3 B4 two SMALL_N near1 _TBL_log.c sin.S sin_return casebase __cos.S constant one pp1 pp2 qq1 qq2 __cos_return q1 q2 q3 q4 __sin.S constant one pp1 pp2 qq1 qq2 __sin_return p1 p2 p3 p4 _TBL_cos.c sccsid _TBL_sin.c sccsid sqrt.S quickreturn constant x y NaN odd two54 insqrt half tmp one twom27 twom57 tfsr nfsr ofsr invalid onehalf onemulp quickcrank table sqrt_return __rem_pio2.S notsmall constant pio2_1 pio2_2 pio2_3 rem_return two24 allarg half pio2_3t pio2_2t pio2_1t zero invpio2 pio2 pio4 medfinal pio2_1t5 finishup _SVID_error.c fmaxx fminx sccsid PI_RZx NaNx setexception Infx matherr.c sccsid _TBL_ipio2.c sccsid __rem_pio2m.c sccsid two24 one zero twon24 init_jk pio2_inf ieee_func.S constant huge scalbn_finite scalbn_return x y two54 scalbn_overflow twom54 tiny scalbn_underflow rndint.S mhalf constant anint_return x irintdata two52 mzero half mtwo52 tmp one zero aint_return rint.S mhalf constant x two52 mzero half mtwo52 tmp one zero rint_return crtn.s __matherr __sqrt __isnormal __cos _SVID_libm_err _start naf_puiss2 nint i_compl_pdivdoubl naf_iniwin _START_ _TBL_cos_hi matherr i_compl_log10 __huge_val _environ _end i_compl_div .stret8 _TBL_log2_lo copysign __expm1 naf_cleannaf _TBL_cos_lo _iob g_NAFVariable i_compl_sub i_compl_log _GLOBAL_OFFSET_TABLE_ cree_list_fenetre_naf i_compl_conj isnormal irint _TBL_ipio2_inf naf_prtabs ilogb isinf atexit exit i_compl_cmplx i_compl_pow i_compl_pow2d i_compl_add log naf_smoy aint i_compl_div2d __copysign malloc rint i_compl_tanh naf_initnaf_notab pow naf_correction i_compl_pmul __log i_compl_div4d __atan2 _init sinh __pow anint fabs .mul __rem_pio2 i_compl_cosh .rem issubnormal i_compl_pmuldoubl signbit __atan naf_four1 naf_mftnaf expm1 sqrt i_compl_exp hypot _END_ _TBL_log_hi i_compl_sinh _DYNAMIC naf_inifre naf_cleannaf_notab printf __iob i_compl_module __signbit i_compl_angle __cosh _TBL_log_lo _TBL_atan_hi naf_initnaf i_compl_powreel _TBL_sin_hi atan2 i_compl_mul __nint _TBL_exp2_hi _exit delete_list_fenetre_naf iszero __iszero exp environ errno _TBL_sin_lo __cg89_used scalbn __exp __scalbn free _TBL_atan_lo _write __irint __rem_pio2m _edata _PROCEDURE_LINKAGE_TABLE_ i_compl_cos __ilogb __isinf _TBL_exp2_lo concat_list_fenetre_naf _etext _lib_version i_compl_psub fflush __aint atan i_compl_pdiv __rint i_compl_sin main pi i_compl_muldoubl .div naf_tessol __sinh __fabs __anint __k_sin _TBL_log2_hi _fini i_compl_paddconst sin __hypot i_compl_padd __issubnormal __k_cos fprintf i_compl_tan cosh __sin cos  @(#)crti.s	1.2	89/12/08 SMI  @(#)crt1.s	1.2	89/12/08 SMI @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI @(#)__fstd.S 1.2 92/05/28 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 20 Aug 1992
 @(#)values-Xt.c	1.6	89/10/24 SMI @(#)synonyms.h	1.5	89/12/18 SMI @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.12 92/04/17 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 20 Aug 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)stdio.h	1.69	98/07/13 SMI @(#)feature_tests.h	1.17	97/12/04 SMI @(#)isa_defs.h	1.15	97/11/22 SMI @(#)va_list.h	1.11	97/11/22 SMI @(#)stdio_tag.h	1.3	98/04/20 SMI @(#)stdio_impl.h	1.7	98/04/17 SMI @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)sunmath.h	1.5	92/04/29 @(#)float.h	1.15	97/11/22 SMI @(#)stdlib.h	1.44	98/01/22 SMI acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)stdio.h	1.69	98/07/13 SMI @(#)feature_tests.h	1.17	97/12/04 SMI @(#)isa_defs.h	1.15	97/11/22 SMI @(#)va_list.h	1.11	97/11/22 SMI @(#)stdio_tag.h	1.3	98/04/20 SMI @(#)stdio_impl.h	1.7	98/04/17 SMI @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)sunmath.h	1.5	92/04/29 @(#)float.h	1.15	97/11/22 SMI @(#)stdlib.h	1.44	98/01/22 SMI acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)errno.h	1.2	90/03/28 SMI @(#)errno.h	1.6	89/11/15 SMI @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)sunmath.h	1.5	92/04/29 @(#)unistd.h	1.2	90/03/30 SMI @(#)types.h	1.5	90/01/05 SMI @(#)machtypes.h	1.3	90/01/20 SMI @(#)select.h	1.4	89/11/09 SMI @(#)time.h	1.2	90/05/11 SMI @(#)time.h	1.2	90/03/30 SMI @(#)unistd.h	1.3	91/12/10 SMI acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)ieeefp.h	1.6 92/04/15 SunPro @(#)math.h	1.75	92/06/23 @(#)floatingpoint.h	1.13 92/08/25 SunPro @(#)stdio.h	1.2	90/03/29 SMI @(#)sunmath.h	1.5	92/04/29 acomp: (CDS) SPARCompilers 2.0.1 03 Sep 1992  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  as: C Development Set  (CDS) SPARCompilers 2.0.1 03 Sep 1992
 @(#)asm_linkage.h	1.10	90/01/08 SMI @(#)stack.h	1.1	91/07/24 SMI @(#)trap.h	1.2	90/09/13 SMI  @(#)crtn.s	1.2	89/12/08 SMI ld: Software Generation Utilities - Solaris/ELF (3.0)             �   d          Gd         g8          �8          \<                z   d          0d         L8          p8          <<          G*                u   d          0d         G8          k8          <<                �   	d          @d         ^8          �8          S<                �   	d          @d         ^8          �8          S<                �   d          >d         Z8          ~8          O<                �   d          Dd         f8          �8          [<                �   d          Dd         f8          �8          [<                �   d          ?d         \8          �8          Q<                �   d          ?d         \8          �8          Q<                �   	d          @d         ^8          �8          S<                �   d          Dd         f8          �8          [<                �   d          Cd         d8          �8          Y<                �   d          Cd         d8          �8          Y<                �   d          Cd         d8          �8          Y<                �   d          Fd         j8          �8          _<                �   d          Bd         b8          �8          W<                �   d          Ed         h8          �8          ]<                �   d          Fd         j8          �8          _<        .interp .hash .dynsym .dynstr .SUNW_version .rela.bss .rela.plt .text .init .fini .rodata .rodata1 .got .plt .dynamic .data .data1 .bss .symtab .strtab .comment .stab.index .shstrtab .stab.indexstr  values-Xt.c /export/set/pergolesi/bootstrap/2.0.1/lang/libansi/sparc/ ../src/values-Xt.c   Xt ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/values-xt.o  example.c /home/pecan1/acct/csteier/simu/naff/ example.c   Xa ; V=2.0 main /home/pecan1/acct/csteier/simu/naff example.o  modnaff.c /home/pecan1/acct/csteier/simu/naff/ modnaff.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff modnaff.o  hypot.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/hypot.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(hypot.o)  atan2.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/atan2.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(atan2.o)  pow.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/pow.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(pow.o)  _TBL_exp2.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_exp2.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_exp2.o)  _TBL_log2.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_log2.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_log2.o)  cosh.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/cosh.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(cosh.o)  sinh.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/sinh.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(sinh.o)  expm1.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/expm1.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(expm1.o)  _TBL_atan.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_atan.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_atan.o)  _TBL_log.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_log.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_log.o)  _TBL_cos.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_cos.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_cos.o)  _TBL_sin.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_sin.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_sin.o)  _SVID_error.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_SVID_error.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_SVID_error.o)  matherr.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/matherr.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(matherr.o)  _TBL_ipio2.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/_TBL_ipio2.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(_TBL_ipio2.o)  __rem_pio2m.c /export/set/pergolesi/bootstrap/2.0.1/lang/libm/sparc/ ../src/C/__rem_pio2m.c   Xa ; V=2.0 /home/pecan1/acct/csteier/simu/naff /opt/SUNWspro-2.0/bin/../SC2.0.1/libm.a(__rem_pio2m.o)                                                      �   �                     	        �   �  $                                                      �                  o���    �  �                    -            $               7       8  8   �               A       �  � )t                  G       GH GH                     M       GT GT                     S       G` G`  1                   [       x` x`  �                  d       � �                    i       � �   �                 n       �� ��   �                w       �� ��  �                  }       �p �p   �                  �       �h �h  �                  �            �h        [         �            ��  .                  �            ��  �                  �            ݬ  d                 �            �   �                  �            ��  C               